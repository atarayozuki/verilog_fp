`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:48:49 06/20/2012 
// Design Name: 
// Module Name:    fp 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module fp(appsel,bck,c4,cs1,cs2,data,db0,db1,db2,db3,db4,db5,db6,db7,di,dl,dn,dr,dt,en,l1,l2,l3,l4,ld,ld0000,ld0001,ld0010,ld0011,ld0100,ld0101,ld0110,ld0111,ld1000,ld1001,ld1010,ld1011,ld1100,ld1101,ld1110,ld1111,lu,md,ml,mr,mu,rd,rst,ru,rw,sysclk,ul,up,ur,ws,clk,d5,d6,d7,d8,r1/*,r2*/,r3,s1,s4/*,s6*/,s8
    );
output appsel,bck,c4,cs1,cs2,data,db0,db1,db2,db3,db4,db5,db6,db7,di,dl,dn,dr,dt,en,l1,l2,l3,l4,ld,ld0000,ld0001,ld0010,ld0011,ld0100,ld0101,ld0110,ld0111,ld1000,ld1001,ld1010,ld1011,ld1100,ld1101,ld1110,ld1111,lu,md,ml,mr,mu,rd,rst,ru,rw,sysclk,ul,up,ur,ws;
input  clk,d5,d6,d7,d8,r1/*,r2*/,r3,s1,s4/*,s6*/,s8;

reg    m0000000_0;
reg    m0000000_1;
reg    m0000001_0;
reg    m0000001_1;
reg    m0000010_0;
reg    m0000010_1;
reg    m0000011_0;
reg    m0000011_1;
reg    m0000100_0;
reg    m0000100_1;
reg    m0000101_0;
reg    m0000101_1;
reg    m0000110_0;
reg    m0000110_1;
reg    m0000111_0;
reg    m0000111_1;
reg    m0001000_0;
reg    m0001000_1;
reg    m0001001_0;
reg    m0001001_1;
reg    m0001010_0;
reg    m0001010_1;
reg    m0001011_0;
reg    m0001011_1;
reg    m0001100_0;
reg    m0001100_1;
reg    m0001101_0;
reg    m0001101_1;
reg    m0001110_0;
reg    m0001110_1;
reg    m0001111_0;
reg    m0001111_1;
reg    m0010000_0;
reg    m0010000_1;
reg    m0010001_0;
reg    m0010001_1;
reg    m0010010_0;
reg    m0010010_1;
reg    m0010011_0;
reg    m0010011_1;
reg    m0010100_0;
reg    m0010100_1;
reg    m0010101_0;
reg    m0010101_1;
reg    m0010110_0;
reg    m0010110_1;
reg    m0010111_0;
reg    m0010111_1;
reg    m0011000_0;
reg    m0011000_1;
reg    m0011001_0;
reg    m0011001_1;
reg    m0011010_0;
reg    m0011010_1;
reg    m0011011_0;
reg    m0011011_1;
reg    m0011100_0;
reg    m0011100_1;
reg    m0011101_0;
reg    m0011101_1;
reg    m0011110_0;
reg    m0011110_1;
reg    m0011111_0;
reg    m0011111_1;
reg    m0100000_0;
reg    m0100000_1;
reg    m0100001_0;
reg    m0100001_1;
reg    m0100010_0;
reg    m0100010_1;
reg    m0100011_0;
reg    m0100011_1;
reg    m0100100_0;
reg    m0100100_1;
reg    m0100101_0;
reg    m0100101_1;
reg    m0100110_0;
reg    m0100110_1;
reg    m0100111_0;
reg    m0100111_1;
reg    m0101000_0;
reg    m0101000_1;
reg    m0101001_0;
reg    m0101001_1;
reg    m0101010_0;
reg    m0101010_1;
reg    m0101011_0;
reg    m0101011_1;
reg    m0101100_0;
reg    m0101100_1;
reg    m0101101_0;
reg    m0101101_1;
reg    m0101110_0;
reg    m0101110_1;
reg    m0101111_0;
reg    m0101111_1;
reg    m0110000_0;
reg    m0110000_1;
reg    m0110001_0;
reg    m0110001_1;
reg    m0110010_0;
reg    m0110010_1;
reg    m0110011_0;
reg    m0110011_1;
reg    m0110100_0;
reg    m0110100_1;
reg    m0110101_0;
reg    m0110101_1;
reg    m0110110_0;
reg    m0110110_1;
reg    m0110111_0;
reg    m0110111_1;
reg    m0111000_0;
reg    m0111000_1;
reg    m0111001_0;
reg    m0111001_1;
reg    m0111010_0;
reg    m0111010_1;
reg    m0111011_0;
reg    m0111011_1;
reg    m0111100_0;
reg    m0111100_1;
reg    m0111101_0;
reg    m0111101_1;
reg    m0111110_0;
reg    m0111110_1;
reg    m0111111_0;
reg    m0111111_1;
reg    m1000000_0;
reg    m1000000_1;
reg    m1000001_0;
reg    m1000001_1;
reg    m1000010_0;
reg    m1000010_1;
reg    m1000011_0;
reg    m1000011_1;
reg    m1000100_0;
reg    m1000100_1;
reg    m1000101_0;
reg    m1000101_1;
reg    m1000110_0;
reg    m1000110_1;
reg    m1000111_0;
reg    m1000111_1;
reg    m1001000_0;
reg    m1001000_1;
reg    m1001001_0;
reg    m1001001_1;
reg    m1001010_0;
reg    m1001010_1;
reg    m1001011_0;
reg    m1001011_1;
reg    m1001100_0;
reg    m1001100_1;
reg    m1001101_0;
reg    m1001101_1;
reg    m1001110_0;
reg    m1001110_1;
reg    m1001111_0;
reg    m1001111_1;
reg    m1010000_0;
reg    m1010000_1;
reg    m1010001_0;
reg    m1010001_1;
reg    m1010010_0;
reg    m1010010_1;
reg    m1010011_0;
reg    m1010011_1;
reg    m1010100_0;
reg    m1010100_1;
reg    m1010101_0;
reg    m1010101_1;
reg    m1010110_0;
reg    m1010110_1;
reg    m1010111_0;
reg    m1010111_1;
reg    m1011000_0;
reg    m1011000_1;
reg    m1011001_0;
reg    m1011001_1;
reg    m1011010_0;
reg    m1011010_1;
reg    m1011011_0;
reg    m1011011_1;
reg    m1011100_0;
reg    m1011100_1;
reg    m1011101_0;
reg    m1011101_1;
reg    m1011110_0;
reg    m1011110_1;
reg    m1011111_0;
reg    m1011111_1;
reg    m1100000_0;
reg    m1100000_1;
reg    m1100001_0;
reg    m1100001_1;
reg    m1100010_0;
reg    m1100010_1;
reg    m1100011_0;
reg    m1100011_1;
reg    m1100100_0;
reg    m1100100_1;
reg    m1100101_0;
reg    m1100101_1;
reg    m1100110_0;
reg    m1100110_1;
reg    m1100111_0;
reg    m1100111_1;
reg    m1101000_0;
reg    m1101000_1;
reg    m1101001_0;
reg    m1101001_1;
reg    m1101010_0;
reg    m1101010_1;
reg    m1101011_0;
reg    m1101011_1;
reg    m1101100_0;
reg    m1101100_1;
reg    m1101101_0;
reg    m1101101_1;
reg    m1101110_0;
reg    m1101110_1;
reg    m1101111_0;
reg    m1101111_1;
reg    m1110000_0;
reg    m1110000_1;
reg    m1110001_0;
reg    m1110001_1;
reg    m1110010_0;
reg    m1110010_1;
reg    m1110011_0;
reg    m1110011_1;
reg    m1110100_0;
reg    m1110100_1;
reg    m1110101_0;
reg    m1110101_1;
reg    m1110110_0;
reg    m1110110_1;
reg    m1110111_0;
reg    m1110111_1;
reg    m1111000_0;
reg    m1111000_1;
reg    m1111001_0;
reg    m1111001_1;
reg    m1111010_0;
reg    m1111010_1;
reg    m1111011_0;
reg    m1111011_1;
reg    m1111100_0;
reg    m1111100_1;
reg    m1111101_0;
reg    m1111101_1;
reg    m1111110_0;
reg    m1111110_1;
reg    m1111111_0;
reg    m1111111_1;

reg    q0000000_0;
reg    q0000000_1;
reg    q0000001_0;
reg    q0000001_1;
reg    q0000010_0;
reg    q0000010_1;
reg    q0000011_0;
reg    q0000011_1;
reg    q0000100_0;
reg    q0000100_1;
reg    q0000101_0;
reg    q0000101_1;
reg    q0000110_0;
reg    q0000110_1;
reg    q0000111_0;
reg    q0000111_1;
reg    q0001000_0;
reg    q0001000_1;
reg    q0001001_0;
reg    q0001001_1;
reg    q0001010_0;
reg    q0001010_1;
reg    q0001011_0;
reg    q0001011_1;
reg    q0001100_0;
reg    q0001100_1;
reg    q0001101_0;
reg    q0001101_1;
reg    q0001110_0;
reg    q0001110_1;
reg    q0001111_0;
reg    q0001111_1;
reg    q0010000_0;
reg    q0010000_1;
reg    q0010001_0;
reg    q0010001_1;
reg    q0010010_0;
reg    q0010010_1;
reg    q0010011_0;
reg    q0010011_1;
reg    q0010100_0;
reg    q0010100_1;
reg    q0010101_0;
reg    q0010101_1;
reg    q0010110_0;
reg    q0010110_1;
reg    q0010111_0;
reg    q0010111_1;
reg    q0011000_0;
reg    q0011000_1;
reg    q0011001_0;
reg    q0011001_1;
reg    q0011010_0;
reg    q0011010_1;
reg    q0011011_0;
reg    q0011011_1;
reg    q0011100_0;
reg    q0011100_1;
reg    q0011101_0;
reg    q0011101_1;
reg    q0011110_0;
reg    q0011110_1;
reg    q0011111_0;
reg    q0011111_1;
reg    q0100000_0;
reg    q0100000_1;
reg    q0100001_0;
reg    q0100001_1;
reg    q0100010_0;
reg    q0100010_1;
reg    q0100011_0;
reg    q0100011_1;
reg    q0100100_0;
reg    q0100100_1;
reg    q0100101_0;
reg    q0100101_1;
reg    q0100110_0;
reg    q0100110_1;
reg    q0100111_0;
reg    q0100111_1;
reg    q0101000_0;
reg    q0101000_1;
reg    q0101001_0;
reg    q0101001_1;
reg    q0101010_0;
reg    q0101010_1;
reg    q0101011_0;
reg    q0101011_1;
reg    q0101100_0;
reg    q0101100_1;
reg    q0101101_0;
reg    q0101101_1;
reg    q0101110_0;
reg    q0101110_1;
reg    q0101111_0;
reg    q0101111_1;
reg    q0110000_0;
reg    q0110000_1;
reg    q0110001_0;
reg    q0110001_1;
reg    q0110010_0;
reg    q0110010_1;
reg    q0110011_0;
reg    q0110011_1;
reg    q0110100_0;
reg    q0110100_1;
reg    q0110101_0;
reg    q0110101_1;
reg    q0110110_0;
reg    q0110110_1;
reg    q0110111_0;
reg    q0110111_1;
reg    q0111000_0;
reg    q0111000_1;
reg    q0111001_0;
reg    q0111001_1;
reg    q0111010_0;
reg    q0111010_1;
reg    q0111011_0;
reg    q0111011_1;
reg    q0111100_0;
reg    q0111100_1;
reg    q0111101_0;
reg    q0111101_1;
reg    q0111110_0;
reg    q0111110_1;
reg    q0111111_0;
reg    q0111111_1;
reg    q1000000_0;
reg    q1000000_1;
reg    q1000001_0;
reg    q1000001_1;
reg    q1000010_0;
reg    q1000010_1;
reg    q1000011_0;
reg    q1000011_1;
reg    q1000100_0;
reg    q1000100_1;
reg    q1000101_0;
reg    q1000101_1;
reg    q1000110_0;
reg    q1000110_1;
reg    q1000111_0;
reg    q1000111_1;
reg    q1001000_0;
reg    q1001000_1;
reg    q1001001_0;
reg    q1001001_1;
reg    q1001010_0;
reg    q1001010_1;
reg    q1001011_0;
reg    q1001011_1;
reg    q1001100_0;
reg    q1001100_1;
reg    q1001101_0;
reg    q1001101_1;
reg    q1001110_0;
reg    q1001110_1;
reg    q1001111_0;
reg    q1001111_1;
reg    q1010000_0;
reg    q1010000_1;
reg    q1010001_0;
reg    q1010001_1;
reg    q1010010_0;
reg    q1010010_1;
reg    q1010011_0;
reg    q1010011_1;
reg    q1010100_0;
reg    q1010100_1;
reg    q1010101_0;
reg    q1010101_1;
reg    q1010110_0;
reg    q1010110_1;
reg    q1010111_0;
reg    q1010111_1;
reg    q1011000_0;
reg    q1011000_1;
reg    q1011001_0;
reg    q1011001_1;
reg    q1011010_0;
reg    q1011010_1;
reg    q1011011_0;
reg    q1011011_1;
reg    q1011100_0;
reg    q1011100_1;
reg    q1011101_0;
reg    q1011101_1;
reg    q1011110_0;
reg    q1011110_1;
reg    q1011111_0;
reg    q1011111_1;
reg    q1100000_0;
reg    q1100000_1;
reg    q1100001_0;
reg    q1100001_1;
reg    q1100010_0;
reg    q1100010_1;
reg    q1100011_0;
reg    q1100011_1;
reg    q1100100_0;
reg    q1100100_1;
reg    q1100101_0;
reg    q1100101_1;
reg    q1100110_0;
reg    q1100110_1;
reg    q1100111_0;
reg    q1100111_1;
reg    q1101000_0;
reg    q1101000_1;
reg    q1101001_0;
reg    q1101001_1;
reg    q1101010_0;
reg    q1101010_1;
reg    q1101011_0;
reg    q1101011_1;
reg    q1101100_0;
reg    q1101100_1;
reg    q1101101_0;
reg    q1101101_1;
reg    q1101110_0;
reg    q1101110_1;
reg    q1101111_0;
reg    q1101111_1;
reg    q1110000_0;
reg    q1110000_1;
reg    q1110001_0;
reg    q1110001_1;
reg    q1110010_0;
reg    q1110010_1;
reg    q1110011_0;
reg    q1110011_1;
reg    q1110100_0;
reg    q1110100_1;
reg    q1110101_0;
reg    q1110101_1;
reg    q1110110_0;
reg    q1110110_1;
reg    q1110111_0;
reg    q1110111_1;
reg    q1111000_0;
reg    q1111000_1;
reg    q1111001_0;
reg    q1111001_1;
reg    q1111010_0;
reg    q1111010_1;
reg    q1111011_0;
reg    q1111011_1;
reg    q1111100_0;
reg    q1111100_1;
reg    q1111101_0;
reg    q1111101_1;
reg    q1111110_0;
reg    q1111110_1;
reg    q1111111_0;
reg    q1111111_1;

reg    m000000_0;
reg    m000000_1;
reg    m000001_0;
reg    m000001_1;
reg    m000010_0;
reg    m000010_1;
reg    m000011_0;
reg    m000011_1;
reg    m000100_0;
reg    m000100_1;
reg    m000101_0;
reg    m000101_1;
reg    m000110_0;
reg    m000110_1;
reg    m000111_0;
reg    m000111_1;
reg    m001000_0;
reg    m001000_1;
reg    m001001_0;
reg    m001001_1;
reg    m001010_0;
reg    m001010_1;
reg    m001011_0;
reg    m001011_1;
reg    m001100_0;
reg    m001100_1;
reg    m001101_0;
reg    m001101_1;
reg    m001110_0;
reg    m001110_1;
reg    m001111_0;
reg    m001111_1;
reg    m010000_0;
reg    m010000_1;
reg    m010001_0;
reg    m010001_1;
reg    m010010_0;
reg    m010010_1;
reg    m010011_0;
reg    m010011_1;
reg    m010100_0;
reg    m010100_1;
reg    m010101_0;
reg    m010101_1;
reg    m010110_0;
reg    m010110_1;
reg    m010111_0;
reg    m010111_1;
reg    m011000_0;
reg    m011000_1;
reg    m011001_0;
reg    m011001_1;
reg    m011010_0;
reg    m011010_1;
reg    m011011_0;
reg    m011011_1;
reg    m011100_0;
reg    m011100_1;
reg    m011101_0;
reg    m011101_1;
reg    m011110_0;
reg    m011110_1;
reg    m011111_0;
reg    m011111_1;
reg    m100000_0;
reg    m100000_1;
reg    m100001_0;
reg    m100001_1;
reg    m100010_0;
reg    m100010_1;
reg    m100011_0;
reg    m100011_1;
reg    m100100_0;
reg    m100100_1;
reg    m100101_0;
reg    m100101_1;
reg    m100110_0;
reg    m100110_1;
reg    m100111_0;
reg    m100111_1;
reg    m101000_0;
reg    m101000_1;
reg    m101001_0;
reg    m101001_1;
reg    m101010_0;
reg    m101010_1;
reg    m101011_0;
reg    m101011_1;
reg    m101100_0;
reg    m101100_1;
reg    m101101_0;
reg    m101101_1;
reg    m101110_0;
reg    m101110_1;
reg    m101111_0;
reg    m101111_1;
reg    m110000_0;
reg    m110000_1;
reg    m110001_0;
reg    m110001_1;
reg    m110010_0;
reg    m110010_1;
reg    m110011_0;
reg    m110011_1;
reg    m110100_0;
reg    m110100_1;
reg    m110101_0;
reg    m110101_1;
reg    m110110_0;
reg    m110110_1;
reg    m110111_0;
reg    m110111_1;
reg    m111000_0;
reg    m111000_1;
reg    m111001_0;
reg    m111001_1;
reg    m111010_0;
reg    m111010_1;
reg    m111011_0;
reg    m111011_1;
reg    m111100_0;
reg    m111100_1;
reg    m111101_0;
reg    m111101_1;
reg    m111110_0;
reg    m111110_1;
reg    m111111_0;
reg    m111111_1;

reg    q000000_0;
reg    q000000_1;
reg    q000001_0;
reg    q000001_1;
reg    q000010_0;
reg    q000010_1;
reg    q000011_0;
reg    q000011_1;
reg    q000100_0;
reg    q000100_1;
reg    q000101_0;
reg    q000101_1;
reg    q000110_0;
reg    q000110_1;
reg    q000111_0;
reg    q000111_1;
reg    q001000_0;
reg    q001000_1;
reg    q001001_0;
reg    q001001_1;
reg    q001010_0;
reg    q001010_1;
reg    q001011_0;
reg    q001011_1;
reg    q001100_0;
reg    q001100_1;
reg    q001101_0;
reg    q001101_1;
reg    q001110_0;
reg    q001110_1;
reg    q001111_0;
reg    q001111_1;
reg    q010000_0;
reg    q010000_1;
reg    q010001_0;
reg    q010001_1;
reg    q010010_0;
reg    q010010_1;
reg    q010011_0;
reg    q010011_1;
reg    q010100_0;
reg    q010100_1;
reg    q010101_0;
reg    q010101_1;
reg    q010110_0;
reg    q010110_1;
reg    q010111_0;
reg    q010111_1;
reg    q011000_0;
reg    q011000_1;
reg    q011001_0;
reg    q011001_1;
reg    q011010_0;
reg    q011010_1;
reg    q011011_0;
reg    q011011_1;
reg    q011100_0;
reg    q011100_1;
reg    q011101_0;
reg    q011101_1;
reg    q011110_0;
reg    q011110_1;
reg    q011111_0;
reg    q011111_1;
reg    q100000_0;
reg    q100000_1;
reg    q100001_0;
reg    q100001_1;
reg    q100010_0;
reg    q100010_1;
reg    q100011_0;
reg    q100011_1;
reg    q100100_0;
reg    q100100_1;
reg    q100101_0;
reg    q100101_1;
reg    q100110_0;
reg    q100110_1;
reg    q100111_0;
reg    q100111_1;
reg    q101000_0;
reg    q101000_1;
reg    q101001_0;
reg    q101001_1;
reg    q101010_0;
reg    q101010_1;
reg    q101011_0;
reg    q101011_1;
reg    q101100_0;
reg    q101100_1;
reg    q101101_0;
reg    q101101_1;
reg    q101110_0;
reg    q101110_1;
reg    q101111_0;
reg    q101111_1;
reg    q110000_0;
reg    q110000_1;
reg    q110001_0;
reg    q110001_1;
reg    q110010_0;
reg    q110010_1;
reg    q110011_0;
reg    q110011_1;
reg    q110100_0;
reg    q110100_1;
reg    q110101_0;
reg    q110101_1;
reg    q110110_0;
reg    q110110_1;
reg    q110111_0;
reg    q110111_1;
reg    q111000_0;
reg    q111000_1;
reg    q111001_0;
reg    q111001_1;
reg    q111010_0;
reg    q111010_1;
reg    q111011_0;
reg    q111011_1;
reg    q111100_0;
reg    q111100_1;
reg    q111101_0;
reg    q111101_1;
reg    q111110_0;
reg    q111110_1;
reg    q111111_0;
reg    q111111_1;

reg    m0001;
reg    m0002;
reg    m0003;
reg    m0004;
reg    m0005;
reg    m0006;
reg    m0007;
reg    m0008;
reg    m0009;
reg    m0010;
reg    m0011;
reg    m0012;
reg    m0013;
reg    m0014;
reg    m0015;
reg    m0016;
reg    m0017;
reg    m0018;
reg    m0019;
reg    m0020;
reg    m0021;
reg    m0022;
reg    m0023;
reg    m0024;
reg    m0025;
reg    m0026;
reg    m0027;
reg    m0028;
reg    m0029;
reg    m0030;

reg    q0001;
reg    q0002;
reg    q0003;
reg    q0004;
reg    q0005;
reg    q0006;
reg    q0007;
reg    q0008;
reg    q0009;
reg    q0010;
reg    q0011;
reg    q0012;
reg    q0013;
reg    q0014;
reg    q0015;
reg    q0016;
reg    q0017;
reg    q0018;
reg    q0019;
reg    q0020;
reg    q0021;
reg    q0022;
reg    q0023;
reg    q0024;
reg    q0025;
reg    q0026;
reg    q0027;
reg    q0028;
reg    q0029;
reg    q0030;
//x
reg    m0031;
reg    m0032;
reg    m0033;
reg    m0034;
reg    m0035;
reg    m0036;
reg    m0037;
reg    m0038;
reg    m0039;
reg    m0040;
reg    m0041;
reg    m0042;
reg    m0043;
reg    m0044;
reg    m0045;
reg    m0046;
reg    m0047;
reg    m0048;
reg    m0049;
reg    m0050;
reg    m0051;
reg    m0052;
reg    m0053;
reg    m0054;
reg    m0055;
reg    m0056;
reg    m0057;
reg    m0058;
reg    m0059;
reg    m0060;

reg    q0031;
reg    q0032;
reg    q0033;
reg    q0034;
reg    q0035;
reg    q0036;
reg    q0037;
reg    q0038;
reg    q0039;
reg    q0040;
reg    q0041;
reg    q0042;
reg    q0043;
reg    q0044;
reg    q0045;
reg    q0046;
reg    q0047;
reg    q0048;
reg    q0049;
reg    q0050;
reg    q0051;
reg    q0052;
reg    q0053;
reg    q0054;
reg    q0055;
reg    q0056;
reg    q0057;
reg    q0058;
reg    q0059;
reg    q0060;

reg    m0061;
reg    m0062;
reg    m0063;
reg    m0064;
reg    m0065;
reg    m0066;
reg    m0067;
reg    m0068;
reg    m0069;
reg    m0070;
reg    m0071;
reg    m0072;
reg    m0073;
reg    m0074;
reg    m0075;
reg    m0076;
reg    m0077;
reg    m0078;
reg    m0079;
reg    m0080;
reg    m0081;
reg    m0082;
reg    m0083;
reg    m0084;
reg    m0085;
reg    m0086;
reg    m0087;
reg    m0088;
reg    m0089;
reg    m0090;

reg    q0061;
reg    q0062;
reg    q0063;
reg    q0064;
reg    q0065;
reg    q0066;
reg    q0067;
reg    q0068;
reg    q0069;
reg    q0070;
reg    q0071;
reg    q0072;
reg    q0073;
reg    q0074;
reg    q0075;
reg    q0076;
reg    q0077;
reg    q0078;
reg    q0079;
reg    q0080;
reg    q0081;
reg    q0082;
reg    q0083;
reg    q0084;
reg    q0085;
reg    q0086;
reg    q0087;
reg    q0088;
reg    q0089;
reg    q0090;
//y
reg    m0091;
reg    m0092;
reg    m0093;
reg    m0094;
reg    m0095;
reg    m0096;
reg    m0097;
reg    m0098;
reg    m0099;
reg    m0100;
reg    m0101;
reg    m0102;
reg    m0103;
reg    m0104;
reg    m0105;
reg    m0106;
reg    m0107;
reg    m0108;
reg    m0109;
reg    m0110;
reg    m0111;
reg    m0112;
reg    m0113;
reg    m0114;
reg    m0115;
reg    m0116;
reg    m0117;
reg    m0118;
reg    m0119;
reg    m0120;

reg    q0091;
reg    q0092;
reg    q0093;
reg    q0094;
reg    q0095;
reg    q0096;
reg    q0097;
reg    q0098;
reg    q0099;
reg    q0100;
reg    q0101;
reg    q0102;
reg    q0103;
reg    q0104;
reg    q0105;
reg    q0106;
reg    q0107;
reg    q0108;
reg    q0109;
reg    q0110;
reg    q0111;
reg    q0112;
reg    q0113;
reg    q0114;
reg    q0115;
reg    q0116;
reg    q0117;
reg    q0118;
reg    q0119;
reg    q0120;

reg    m0121;
reg    m0122;
reg    m0123;
reg    m0124;
reg    m0125;
reg    m0126;
reg    m0127;
reg    m0128;
reg    m0129;
reg    m0130;
reg    m0131;
reg    m0132;
reg    m0133;
reg    m0134;
reg    m0135;
reg    m0136;
reg    m0137;
reg    m0138;
reg    m0139;
reg    m0140;
reg    m0141;
reg    m0142;
reg    m0143;
reg    m0144;
reg    m0145;
reg    m0146;
reg    m0147;
reg    m0148;
reg    m0149;
reg    m0150;

reg    q0121;
reg    q0122;
reg    q0123;
reg    q0124;
reg    q0125;
reg    q0126;
reg    q0127;
reg    q0128;
reg    q0129;
reg    q0130;
reg    q0131;
reg    q0132;
reg    q0133;
reg    q0134;
reg    q0135;
reg    q0136;
reg    q0137;
reg    q0138;
reg    q0139;
reg    q0140;
reg    q0141;
reg    q0142;
reg    q0143;
reg    q0144;
reg    q0145;
reg    q0146;
reg    q0147;
reg    q0148;
reg    q0149;
reg    q0150;
//1
reg    m0151;
reg    m0152;
reg    m0153;
reg    m0154;
reg    m0155;
reg    m0156;
reg    m0157;
reg    m0158;
reg    m0159;
reg    m0160;
reg    m0161;
reg    m0162;
reg    m0163;
reg    m0164;
reg    m0165;
reg    m0166;
reg    m0167;
reg    m0168;
reg    m0169;
reg    m0170;
reg    m0171;
reg    m0172;
reg    m0173;
reg    m0174;
reg    m0175;
reg    m0176;
reg    m0177;
reg    m0178;
reg    m0179;
reg    m0180;

reg    q0151;
reg    q0152;
reg    q0153;
reg    q0154;
reg    q0155;
reg    q0156;
reg    q0157;
reg    q0158;
reg    q0159;
reg    q0160;
reg    q0161;
reg    q0162;
reg    q0163;
reg    q0164;
reg    q0165;
reg    q0166;
reg    q0167;
reg    q0168;
reg    q0169;
reg    q0170;
reg    q0171;
reg    q0172;
reg    q0173;
reg    q0174;
reg    q0175;
reg    q0176;
reg    q0177;
reg    q0178;
reg    q0179;
reg    q0180;

reg    m0181;
reg    m0182;
reg    m0183;
reg    m0184;
reg    m0185;
reg    m0186;
reg    m0187;
reg    m0188;
reg    m0189;
reg    m0190;
reg    m0191;
reg    m0192;
reg    m0193;
reg    m0194;
reg    m0195;
reg    m0196;
reg    m0197;
reg    m0198;
reg    m0199;
reg    m0200;
reg    m0201;
reg    m0202;
reg    m0203;
reg    m0204;
reg    m0205;
reg    m0206;
reg    m0207;
reg    m0208;
reg    m0209;
reg    m0210;

reg    q0181;
reg    q0182;
reg    q0183;
reg    q0184;
reg    q0185;
reg    q0186;
reg    q0187;
reg    q0188;
reg    q0189;
reg    q0190;
reg    q0191;
reg    q0192;
reg    q0193;
reg    q0194;
reg    q0195;
reg    q0196;
reg    q0197;
reg    q0198;
reg    q0199;
reg    q0200;
reg    q0201;
reg    q0202;
reg    q0203;
reg    q0204;
reg    q0205;
reg    q0206;
reg    q0207;
reg    q0208;
reg    q0209;
reg    q0210;
//2
reg    m0211;
reg    m0212;
reg    m0213;
reg    m0214;
reg    m0215;
reg    m0216;
reg    m0217;
reg    m0218;
reg    m0219;
reg    m0220;
reg    m0221;
reg    m0222;
reg    m0223;
reg    m0224;
reg    m0225;
reg    m0226;
reg    m0227;
reg    m0228;
reg    m0229;
reg    m0230;
reg    m0231;
reg    m0232;
reg    m0233;
reg    m0234;
reg    m0235;
reg    m0236;
reg    m0237;
reg    m0238;
reg    m0239;
reg    m0240;

reg    q0211;
reg    q0212;
reg    q0213;
reg    q0214;
reg    q0215;
reg    q0216;
reg    q0217;
reg    q0218;
reg    q0219;
reg    q0220;
reg    q0221;
reg    q0222;
reg    q0223;
reg    q0224;
reg    q0225;
reg    q0226;
reg    q0227;
reg    q0228;
reg    q0229;
reg    q0230;
reg    q0231;
reg    q0232;
reg    q0233;
reg    q0234;
reg    q0235;
reg    q0236;
reg    q0237;
reg    q0238;
reg    q0239;
reg    q0240;

reg    m0241;
reg    m0242;
reg    m0243;
reg    m0244;
reg    m0245;
reg    m0246;
reg    m0247;
reg    m0248;
reg    m0249;
reg    m0250;
reg    m0251;
reg    m0252;
reg    m0253;
reg    m0254;
reg    m0255;
reg    m0256;
reg    m0257;
reg    m0258;
reg    m0259;
reg    m0260;
reg    m0261;
reg    m0262;
reg    m0263;
reg    m0264;
reg    m0265;
reg    m0266;
reg    m0267;
reg    m0268;
reg    m0269;
reg    m0270;

reg    q0241;
reg    q0242;
reg    q0243;
reg    q0244;
reg    q0245;
reg    q0246;
reg    q0247;
reg    q0248;
reg    q0249;
reg    q0250;
reg    q0251;
reg    q0252;
reg    q0253;
reg    q0254;
reg    q0255;
reg    q0256;
reg    q0257;
reg    q0258;
reg    q0259;
reg    q0260;
reg    q0261;
reg    q0262;
reg    q0263;
reg    q0264;
reg    q0265;
reg    q0266;
reg    q0267;
reg    q0268;
reg    q0269;
reg    q0270;
//s
reg    m0271;
reg    m0272;
reg    m0273;
reg    m0274;
reg    m0275;
reg    m0276;
reg    m0277;
reg    m0278;
reg    m0279;
reg    m0280;
reg    m0281;
reg    m0282;
reg    m0283;
reg    m0284;
reg    m0285;
reg    m0286;
reg    m0287;
reg    m0288;
reg    m0289;
reg    m0290;
reg    m0291;
reg    m0292;
reg    m0293;
reg    m0294;
reg    m0295;
reg    m0296;
reg    m0297;
reg    m0298;
reg    m0299;
reg    m0300;

reg    q0271;
reg    q0272;
reg    q0273;
reg    q0274;
reg    q0275;
reg    q0276;
reg    q0277;
reg    q0278;
reg    q0279;
reg    q0280;
reg    q0281;
reg    q0282;
reg    q0283;
reg    q0284;
reg    q0285;
reg    q0286;
reg    q0287;
reg    q0288;
reg    q0289;
reg    q0290;
reg    q0291;
reg    q0292;
reg    q0293;
reg    q0294;
reg    q0295;
reg    q0296;
reg    q0297;
reg    q0298;
reg    q0299;
reg    q0300;

reg    m0301;
reg    m0302;
reg    m0303;
reg    m0304;
reg    m0305;
reg    m0306;
reg    m0307;
reg    m0308;
reg    m0309;
reg    m0310;
reg    m0311;
reg    m0312;
reg    m0313;
reg    m0314;
reg    m0315;
reg    m0316;
reg    m0317;
reg    m0318;
reg    m0319;
reg    m0320;
reg    m0321;
reg    m0322;
reg    m0323;
reg    m0324;
reg    m0325;
reg    m0326;
reg    m0327;
reg    m0328;
reg    m0329;
reg    m0330;

reg    q0301;
reg    q0302;
reg    q0303;
reg    q0304;
reg    q0305;
reg    q0306;
reg    q0307;
reg    q0308;
reg    q0309;
reg    q0310;
reg    q0311;
reg    q0312;
reg    q0313;
reg    q0314;
reg    q0315;
reg    q0316;
reg    q0317;
reg    q0318;
reg    q0319;
reg    q0320;
reg    q0321;
reg    q0322;
reg    q0323;
reg    q0324;
reg    q0325;
reg    q0326;
reg    q0327;
reg    q0328;
reg    q0329;
reg    q0330;
//so
reg    m0331;
reg    m0332;
reg    m0333;
reg    m0334;
reg    m0335;
reg    m0336;
reg    m0337;
reg    m0338;
reg    m0339;
reg    m0340;
reg    m0341;
reg    m0342;
reg    m0343;
reg    m0344;
reg    m0345;
reg    m0346;
reg    m0347;
reg    m0348;
reg    m0349;
reg    m0350;
reg    m0351;
reg    m0352;
reg    m0353;
reg    m0354;
reg    m0355;
reg    m0356;
reg    m0357;
reg    m0358;
reg    m0359;
reg    m0360;

reg    q0331;
reg    q0332;
reg    q0333;
reg    q0334;
reg    q0335;
reg    q0336;
reg    q0337;
reg    q0338;
reg    q0339;
reg    q0340;
reg    q0341;
reg    q0342;
reg    q0343;
reg    q0344;
reg    q0345;
reg    q0346;
reg    q0347;
reg    q0348;
reg    q0349;
reg    q0350;
reg    q0351;
reg    q0352;
reg    q0353;
reg    q0354;
reg    q0355;
reg    q0356;
reg    q0357;
reg    q0358;
reg    q0359;
reg    q0360;

reg    m0361;
reg    m0362;
reg    m0363;
reg    m0364;
reg    m0365;
reg    m0366;
reg    m0367;
reg    m0368;
reg    m0369;
reg    m0370;
reg    m0371;
reg    m0372;
reg    m0373;
reg    m0374;
reg    m0375;
reg    m0376;
reg    m0377;
reg    m0378;
reg    m0379;
reg    m0380;
reg    m0381;
reg    m0382;
reg    m0383;
reg    m0384;
reg    m0385;
reg    m0386;
reg    m0387;
reg    m0388;
reg    m0389;
reg    m0390;

reg    q0361;
reg    q0362;
reg    q0363;
reg    q0364;
reg    q0365;
reg    q0366;
reg    q0367;
reg    q0368;
reg    q0369;
reg    q0370;
reg    q0371;
reg    q0372;
reg    q0373;
reg    q0374;
reg    q0375;
reg    q0376;
reg    q0377;
reg    q0378;
reg    q0379;
reg    q0380;
reg    q0381;
reg    q0382;
reg    q0383;
reg    q0384;
reg    q0385;
reg    q0386;
reg    q0387;
reg    q0388;
reg    q0389;
reg    q0390;

reg    m100_0;
reg    m100_1;
reg    m101_0;
reg    m101_1;
reg    m162_0;
reg    m162_1;
reg    m163_0;
reg    m163_1;

reg    q100_0;
reg    q100_1;
reg    q101_0;
reg    q101_1;
reg    q162_0;
reg    q162_1;
reg    q163_0;
reg    q163_1;

reg    m200_0;
reg    m200_1;
reg    m201_0;
reg    m201_1;
reg    m262_0;
reg    m262_1;
reg    m263_0;
reg    m263_1;

reg    q200_0;
reg    q200_1;
reg    q201_0;
reg    q201_1;
reg    q262_0;
reg    q262_1;
reg    q263_0;
reg    q263_1;

reg    m102_0;
reg    m102_1;
reg    m103_0;
reg    m103_1;
reg    m104_0;
reg    m104_1;
reg    m105_0;
reg    m105_1;
reg    m106_0;
reg    m106_1;
reg    m107_0;
reg    m107_1;
reg    m108_0;
reg    m108_1;
reg    m109_0;
reg    m109_1;
reg    m110_0;
reg    m110_1;
reg    m111_0;
reg    m111_1;
reg    m112_0;
reg    m112_1;
reg    m113_0;
reg    m113_1;
reg    m114_0;
reg    m114_1;
reg    m115_0;
reg    m115_1;
reg    m116_0;
reg    m116_1;
reg    m117_0;
reg    m117_1;
reg    m118_0;
reg    m118_1;
reg    m119_0;
reg    m119_1;
reg    m120_0;
reg    m120_1;
reg    m121_0;
reg    m121_1;
reg    m122_0;
reg    m122_1;
reg    m123_0;
reg    m123_1;
reg    m124_0;
reg    m124_1;
reg    m125_0;
reg    m125_1;
reg    m126_0;
reg    m126_1;
reg    m127_0;
reg    m127_1;
reg    m128_0;
reg    m128_1;
reg    m129_0;
reg    m129_1;
reg    m130_0;
reg    m130_1;
reg    m131_0;
reg    m131_1;
reg    m132_0;
reg    m132_1;
reg    m133_0;
reg    m133_1;
reg    m134_0;
reg    m134_1;
reg    m135_0;
reg    m135_1;
reg    m136_0;
reg    m136_1;
reg    m137_0;
reg    m137_1;
reg    m138_0;
reg    m138_1;
reg    m139_0;
reg    m139_1;
reg    m140_0;
reg    m140_1;
reg    m141_0;
reg    m141_1;
reg    m142_0;
reg    m142_1;
reg    m143_0;
reg    m143_1;
reg    m144_0;
reg    m144_1;
reg    m145_0;
reg    m145_1;
reg    m146_0;
reg    m146_1;
reg    m147_0;
reg    m147_1;
reg    m148_0;
reg    m148_1;
reg    m149_0;
reg    m149_1;
reg    m150_0;
reg    m150_1;
reg    m151_0;
reg    m151_1;
reg    m152_0;
reg    m152_1;
reg    m153_0;
reg    m153_1;
reg    m154_0;
reg    m154_1;
reg    m155_0;
reg    m155_1;
reg    m156_0;
reg    m156_1;
reg    m157_0;
reg    m157_1;
reg    m158_0;
reg    m158_1;
reg    m159_0;
reg    m159_1;
reg    m160_0;
reg    m160_1;
reg    m161_0;
reg    m161_1;

reg    q102_0;
reg    q102_1;
reg    q103_0;
reg    q103_1;
reg    q104_0;
reg    q104_1;
reg    q105_0;
reg    q105_1;
reg    q106_0;
reg    q106_1;
reg    q107_0;
reg    q107_1;
reg    q108_0;
reg    q108_1;
reg    q109_0;
reg    q109_1;
reg    q110_0;
reg    q110_1;
reg    q111_0;
reg    q111_1;
reg    q112_0;
reg    q112_1;
reg    q113_0;
reg    q113_1;
reg    q114_0;
reg    q114_1;
reg    q115_0;
reg    q115_1;
reg    q116_0;
reg    q116_1;
reg    q117_0;
reg    q117_1;
reg    q118_0;
reg    q118_1;
reg    q119_0;
reg    q119_1;
reg    q120_0;
reg    q120_1;
reg    q121_0;
reg    q121_1;
reg    q122_0;
reg    q122_1;
reg    q123_0;
reg    q123_1;
reg    q124_0;
reg    q124_1;
reg    q125_0;
reg    q125_1;
reg    q126_0;
reg    q126_1;
reg    q127_0;
reg    q127_1;
reg    q128_0;
reg    q128_1;
reg    q129_0;
reg    q129_1;
reg    q130_0;
reg    q130_1;
reg    q131_0;
reg    q131_1;
reg    q132_0;
reg    q132_1;
reg    q133_0;
reg    q133_1;
reg    q134_0;
reg    q134_1;
reg    q135_0;
reg    q135_1;
reg    q136_0;
reg    q136_1;
reg    q137_0;
reg    q137_1;
reg    q138_0;
reg    q138_1;
reg    q139_0;
reg    q139_1;
reg    q140_0;
reg    q140_1;
reg    q141_0;
reg    q141_1;
reg    q142_0;
reg    q142_1;
reg    q143_0;
reg    q143_1;
reg    q144_0;
reg    q144_1;
reg    q145_0;
reg    q145_1;
reg    q146_0;
reg    q146_1;
reg    q147_0;
reg    q147_1;
reg    q148_0;
reg    q148_1;
reg    q149_0;
reg    q149_1;
reg    q150_0;
reg    q150_1;
reg    q151_0;
reg    q151_1;
reg    q152_0;
reg    q152_1;
reg    q153_0;
reg    q153_1;
reg    q154_0;
reg    q154_1;
reg    q155_0;
reg    q155_1;
reg    q156_0;
reg    q156_1;
reg    q157_0;
reg    q157_1;
reg    q158_0;
reg    q158_1;
reg    q159_0;
reg    q159_1;
reg    q160_0;
reg    q160_1;
reg    q161_0;
reg    q161_1;

reg    m202_0;
reg    m202_1;
reg    m203_0;
reg    m203_1;
reg    m204_0;
reg    m204_1;
reg    m205_0;
reg    m205_1;
reg    m206_0;
reg    m206_1;
reg    m207_0;
reg    m207_1;
reg    m208_0;
reg    m208_1;
reg    m209_0;
reg    m209_1;
reg    m210_0;
reg    m210_1;
reg    m211_0;
reg    m211_1;
reg    m212_0;
reg    m212_1;
reg    m213_0;
reg    m213_1;
reg    m214_0;
reg    m214_1;
reg    m215_0;
reg    m215_1;
reg    m216_0;
reg    m216_1;
reg    m217_0;
reg    m217_1;
reg    m218_0;
reg    m218_1;
reg    m219_0;
reg    m219_1;
reg    m220_0;
reg    m220_1;
reg    m221_0;
reg    m221_1;
reg    m222_0;
reg    m222_1;
reg    m223_0;
reg    m223_1;
reg    m224_0;
reg    m224_1;
reg    m225_0;
reg    m225_1;
reg    m226_0;
reg    m226_1;
reg    m227_0;
reg    m227_1;
reg    m228_0;
reg    m228_1;
reg    m229_0;
reg    m229_1;
reg    m230_0;
reg    m230_1;
reg    m231_0;
reg    m231_1;
reg    m232_0;
reg    m232_1;
reg    m233_0;
reg    m233_1;
reg    m234_0;
reg    m234_1;
reg    m235_0;
reg    m235_1;
reg    m236_0;
reg    m236_1;
reg    m237_0;
reg    m237_1;
reg    m238_0;
reg    m238_1;
reg    m239_0;
reg    m239_1;
reg    m240_0;
reg    m240_1;
reg    m241_0;
reg    m241_1;
reg    m242_0;
reg    m242_1;
reg    m243_0;
reg    m243_1;
reg    m244_0;
reg    m244_1;
reg    m245_0;
reg    m245_1;
reg    m246_0;
reg    m246_1;
reg    m247_0;
reg    m247_1;
reg    m248_0;
reg    m248_1;
reg    m249_0;
reg    m249_1;
reg    m250_0;
reg    m250_1;
reg    m251_0;
reg    m251_1;
reg    m252_0;
reg    m252_1;
reg    m253_0;
reg    m253_1;
reg    m254_0;
reg    m254_1;
reg    m255_0;
reg    m255_1;
reg    m256_0;
reg    m256_1;
reg    m257_0;
reg    m257_1;
reg    m258_0;
reg    m258_1;
reg    m259_0;
reg    m259_1;
reg    m260_0;
reg    m260_1;
reg    m261_0;
reg    m261_1;

reg    q202_0;
reg    q202_1;
reg    q203_0;
reg    q203_1;
reg    q204_0;
reg    q204_1;
reg    q205_0;
reg    q205_1;
reg    q206_0;
reg    q206_1;
reg    q207_0;
reg    q207_1;
reg    q208_0;
reg    q208_1;
reg    q209_0;
reg    q209_1;
reg    q210_0;
reg    q210_1;
reg    q211_0;
reg    q211_1;
reg    q212_0;
reg    q212_1;
reg    q213_0;
reg    q213_1;
reg    q214_0;
reg    q214_1;
reg    q215_0;
reg    q215_1;
reg    q216_0;
reg    q216_1;
reg    q217_0;
reg    q217_1;
reg    q218_0;
reg    q218_1;
reg    q219_0;
reg    q219_1;
reg    q220_0;
reg    q220_1;
reg    q221_0;
reg    q221_1;
reg    q222_0;
reg    q222_1;
reg    q223_0;
reg    q223_1;
reg    q224_0;
reg    q224_1;
reg    q225_0;
reg    q225_1;
reg    q226_0;
reg    q226_1;
reg    q227_0;
reg    q227_1;
reg    q228_0;
reg    q228_1;
reg    q229_0;
reg    q229_1;
reg    q230_0;
reg    q230_1;
reg    q231_0;
reg    q231_1;
reg    q232_0;
reg    q232_1;
reg    q233_0;
reg    q233_1;
reg    q234_0;
reg    q234_1;
reg    q235_0;
reg    q235_1;
reg    q236_0;
reg    q236_1;
reg    q237_0;
reg    q237_1;
reg    q238_0;
reg    q238_1;
reg    q239_0;
reg    q239_1;
reg    q240_0;
reg    q240_1;
reg    q241_0;
reg    q241_1;
reg    q242_0;
reg    q242_1;
reg    q243_0;
reg    q243_1;
reg    q244_0;
reg    q244_1;
reg    q245_0;
reg    q245_1;
reg    q246_0;
reg    q246_1;
reg    q247_0;
reg    q247_1;
reg    q248_0;
reg    q248_1;
reg    q249_0;
reg    q249_1;
reg    q250_0;
reg    q250_1;
reg    q251_0;
reg    q251_1;
reg    q252_0;
reg    q252_1;
reg    q253_0;
reg    q253_1;
reg    q254_0;
reg    q254_1;
reg    q255_0;
reg    q255_1;
reg    q256_0;
reg    q256_1;
reg    q257_0;
reg    q257_1;
reg    q258_0;
reg    q258_1;
reg    q259_0;
reg    q259_1;
reg    q260_0;
reg    q260_1;
reg    q261_0;
reg    q261_1;
/*
reg    m1000_0;
reg    m1000_1;
reg    m1001_0;
reg    m1001_1;
reg    m1010_0;
reg    m1010_1;
reg    m1011_0;
reg    m1011_1;
reg    m1100_0;
reg    m1100_1;
reg    m1101_0;
reg    m1101_1;
reg    m1110_0;
reg    m1110_1;
reg    m1111_0;
reg    m1111_1;

reg    q1000_0;
reg    q1000_1;
reg    q1001_0;
reg    q1001_1;
reg    q1010_0;
reg    q1010_1;
reg    q1011_0;
reg    q1011_1;
reg    q1100_0;
reg    q1100_1;
reg    q1101_0;
reg    q1101_1;
reg    q1110_0;
reg    q1110_1;
reg    q1111_0;
reg    q1111_1;

reg    m2000_0;
reg    m2000_1;
reg    m2001_0;
reg    m2001_1;
reg    m2010_0;
reg    m2010_1;
reg    m2011_0;
reg    m2011_1;
reg    m2100_0;
reg    m2100_1;
reg    m2101_0;
reg    m2101_1;
reg    m2110_0;
reg    m2110_1;
reg    m2111_0;
reg    m2111_1;

reg    q2000_0;
reg    q2000_1;
reg    q2001_0;
reg    q2001_1;
reg    q2010_0;
reg    q2010_1;
reg    q2011_0;
reg    q2011_1;
reg    q2100_0;
reg    q2100_1;
reg    q2101_0;
reg    q2101_1;
reg    q2110_0;
reg    q2110_1;
reg    q2111_0;
reg    q2111_1;
*/
reg    m00_0;
reg    m00_1;
reg    m01_0;
reg    m01_1;
reg    m10_0;
reg    m10_1;
reg    m11_0;
reg    m11_1;

reg    q00_0;
reg    q00_1;
reg    q01_0;
reg    q01_1;
reg    q10_0;
reg    q10_1;
reg    q11_0;
reg    q11_1;

reg    ms_0;
reg    ms_1;

reg    qs_0;
reg    qs_1;

reg    mso_0;
reg    mso_1;

reg    qso_0;
reg    qso_1;

reg    m29_0;
reg    m29_1;
reg    m30_0;
reg    m30_1;
reg    m31_0;
reg    m31_1;
reg    m32_0;
reg    m32_1;
reg    m33_0;
reg    m33_1;
reg    m34_0;
reg    m34_1;
reg    m35_0;
reg    m35_1;
reg    m36_0;
reg    m36_1;
reg    m37_0;
reg    m37_1;
reg    m38_0;
reg    m38_1;
reg    m39_0;
reg    m39_1;
reg    m40_0;
reg    m40_1;
reg    m41_0;
reg    m41_1;
reg    m42_0;
reg    m42_1;
reg    m43_0;
reg    m43_1;
reg    m44_0;
reg    m44_1;
reg    m45_0;
reg    m45_1;
reg    m46_0;
reg    m46_1;
reg    m47_0;
reg    m47_1;
reg    m48_0;
reg    m48_1;
reg    m49_0;
reg    m49_1;
reg    m50_0;
reg    m50_1;

reg    q29_0;
reg    q29_1;
reg    q30_0;
reg    q30_1;
reg    q31_0;
reg    q31_1;
reg    q32_0;
reg    q32_1;
reg    q33_0;
reg    q33_1;
reg    q34_0;
reg    q34_1;
reg    q35_0;
reg    q35_1;
reg    q36_0;
reg    q36_1;
reg    q37_0;
reg    q37_1;
reg    q38_0;
reg    q38_1;
reg    q39_0;
reg    q39_1;
reg    q40_0;
reg    q40_1;
reg    q41_0;
reg    q41_1;
reg    q42_0;
reg    q42_1;
reg    q43_0;
reg    q43_1;
reg    q44_0;
reg    q44_1;
reg    q45_0;
reg    q45_1;
reg    q46_0;
reg    q46_1;
reg    q47_0;
reg    q47_1;
reg    q48_0;
reg    q48_1;
reg    q49_0;
reg    q49_1;
reg    q50_0;
reg    q50_1;

reg    m0_0;/*
reg    m0_1;*/
reg    m1_0;/*
reg    m1_1;*/

reg    q0_0;/*
reg    q0_1;*/
reg    q1_0;/*
reg    q1_1;*/

always @(posedge clk)
m0000000_0<=h0000000_0;
always @(posedge clk)
m0000000_1<=h0000000_1;
always @(posedge clk)
m0000001_0<=h0000001_0;
always @(posedge clk)
m0000001_1<=h0000001_1;
always @(posedge clk)
m0000010_0<=h0000010_0;
always @(posedge clk)
m0000010_1<=h0000010_1;
always @(posedge clk)
m0000011_0<=h0000011_0;
always @(posedge clk)
m0000011_1<=h0000011_1;
always @(posedge clk)
m0000100_0<=h0000100_0;
always @(posedge clk)
m0000100_1<=h0000100_1;
always @(posedge clk)
m0000101_0<=h0000101_0;
always @(posedge clk)
m0000101_1<=h0000101_1;
always @(posedge clk)
m0000110_0<=h0000110_0;
always @(posedge clk)
m0000110_1<=h0000110_1;
always @(posedge clk)
m0000111_0<=h0000111_0;
always @(posedge clk)
m0000111_1<=h0000111_1;
always @(posedge clk)
m0001000_0<=h0001000_0;
always @(posedge clk)
m0001000_1<=h0001000_1;
always @(posedge clk)
m0001001_0<=h0001001_0;
always @(posedge clk)
m0001001_1<=h0001001_1;
always @(posedge clk)
m0001010_0<=h0001010_0;
always @(posedge clk)
m0001010_1<=h0001010_1;
always @(posedge clk)
m0001011_0<=h0001011_0;
always @(posedge clk)
m0001011_1<=h0001011_1;
always @(posedge clk)
m0001100_0<=h0001100_0;
always @(posedge clk)
m0001100_1<=h0001100_1;
always @(posedge clk)
m0001101_0<=h0001101_0;
always @(posedge clk)
m0001101_1<=h0001101_1;
always @(posedge clk)
m0001110_0<=h0001110_0;
always @(posedge clk)
m0001110_1<=h0001110_1;
always @(posedge clk)
m0001111_0<=h0001111_0;
always @(posedge clk)
m0001111_1<=h0001111_1;
always @(posedge clk)
m0010000_0<=h0010000_0;
always @(posedge clk)
m0010000_1<=h0010000_1;
always @(posedge clk)
m0010001_0<=h0010001_0;
always @(posedge clk)
m0010001_1<=h0010001_1;
always @(posedge clk)
m0010010_0<=h0010010_0;
always @(posedge clk)
m0010010_1<=h0010010_1;
always @(posedge clk)
m0010011_0<=h0010011_0;
always @(posedge clk)
m0010011_1<=h0010011_1;
always @(posedge clk)
m0010100_0<=h0010100_0;
always @(posedge clk)
m0010100_1<=h0010100_1;
always @(posedge clk)
m0010101_0<=h0010101_0;
always @(posedge clk)
m0010101_1<=h0010101_1;
always @(posedge clk)
m0010110_0<=h0010110_0;
always @(posedge clk)
m0010110_1<=h0010110_1;
always @(posedge clk)
m0010111_0<=h0010111_0;
always @(posedge clk)
m0010111_1<=h0010111_1;
always @(posedge clk)
m0011000_0<=h0011000_0;
always @(posedge clk)
m0011000_1<=h0011000_1;
always @(posedge clk)
m0011001_0<=h0011001_0;
always @(posedge clk)
m0011001_1<=h0011001_1;
always @(posedge clk)
m0011010_0<=h0011010_0;
always @(posedge clk)
m0011010_1<=h0011010_1;
always @(posedge clk)
m0011011_0<=h0011011_0;
always @(posedge clk)
m0011011_1<=h0011011_1;
always @(posedge clk)
m0011100_0<=h0011100_0;
always @(posedge clk)
m0011100_1<=h0011100_1;
always @(posedge clk)
m0011101_0<=h0011101_0;
always @(posedge clk)
m0011101_1<=h0011101_1;
always @(posedge clk)
m0011110_0<=h0011110_0;
always @(posedge clk)
m0011110_1<=h0011110_1;
always @(posedge clk)
m0011111_0<=h0011111_0;
always @(posedge clk)
m0011111_1<=h0011111_1;
always @(posedge clk)
m0100000_0<=h0100000_0;
always @(posedge clk)
m0100000_1<=h0100000_1;
always @(posedge clk)
m0100001_0<=h0100001_0;
always @(posedge clk)
m0100001_1<=h0100001_1;
always @(posedge clk)
m0100010_0<=h0100010_0;
always @(posedge clk)
m0100010_1<=h0100010_1;
always @(posedge clk)
m0100011_0<=h0100011_0;
always @(posedge clk)
m0100011_1<=h0100011_1;
always @(posedge clk)
m0100100_0<=h0100100_0;
always @(posedge clk)
m0100100_1<=h0100100_1;
always @(posedge clk)
m0100101_0<=h0100101_0;
always @(posedge clk)
m0100101_1<=h0100101_1;
always @(posedge clk)
m0100110_0<=h0100110_0;
always @(posedge clk)
m0100110_1<=h0100110_1;
always @(posedge clk)
m0100111_0<=h0100111_0;
always @(posedge clk)
m0100111_1<=h0100111_1;
always @(posedge clk)
m0101000_0<=h0101000_0;
always @(posedge clk)
m0101000_1<=h0101000_1;
always @(posedge clk)
m0101001_0<=h0101001_0;
always @(posedge clk)
m0101001_1<=h0101001_1;
always @(posedge clk)
m0101010_0<=h0101010_0;
always @(posedge clk)
m0101010_1<=h0101010_1;
always @(posedge clk)
m0101011_0<=h0101011_0;
always @(posedge clk)
m0101011_1<=h0101011_1;
always @(posedge clk)
m0101100_0<=h0101100_0;
always @(posedge clk)
m0101100_1<=h0101100_1;
always @(posedge clk)
m0101101_0<=h0101101_0;
always @(posedge clk)
m0101101_1<=h0101101_1;
always @(posedge clk)
m0101110_0<=h0101110_0;
always @(posedge clk)
m0101110_1<=h0101110_1;
always @(posedge clk)
m0101111_0<=h0101111_0;
always @(posedge clk)
m0101111_1<=h0101111_1;
always @(posedge clk)
m0110000_0<=h0110000_0;
always @(posedge clk)
m0110000_1<=h0110000_1;
always @(posedge clk)
m0110001_0<=h0110001_0;
always @(posedge clk)
m0110001_1<=h0110001_1;
always @(posedge clk)
m0110010_0<=h0110010_0;
always @(posedge clk)
m0110010_1<=h0110010_1;
always @(posedge clk)
m0110011_0<=h0110011_0;
always @(posedge clk)
m0110011_1<=h0110011_1;
always @(posedge clk)
m0110100_0<=h0110100_0;
always @(posedge clk)
m0110100_1<=h0110100_1;
always @(posedge clk)
m0110101_0<=h0110101_0;
always @(posedge clk)
m0110101_1<=h0110101_1;
always @(posedge clk)
m0110110_0<=h0110110_0;
always @(posedge clk)
m0110110_1<=h0110110_1;
always @(posedge clk)
m0110111_0<=h0110111_0;
always @(posedge clk)
m0110111_1<=h0110111_1;
always @(posedge clk)
m0111000_0<=h0111000_0;
always @(posedge clk)
m0111000_1<=h0111000_1;
always @(posedge clk)
m0111001_0<=h0111001_0;
always @(posedge clk)
m0111001_1<=h0111001_1;
always @(posedge clk)
m0111010_0<=h0111010_0;
always @(posedge clk)
m0111010_1<=h0111010_1;
always @(posedge clk)
m0111011_0<=h0111011_0;
always @(posedge clk)
m0111011_1<=h0111011_1;
always @(posedge clk)
m0111100_0<=h0111100_0;
always @(posedge clk)
m0111100_1<=h0111100_1;
always @(posedge clk)
m0111101_0<=h0111101_0;
always @(posedge clk)
m0111101_1<=h0111101_1;
always @(posedge clk)
m0111110_0<=h0111110_0;
always @(posedge clk)
m0111110_1<=h0111110_1;
always @(posedge clk)
m0111111_0<=h0111111_0;
always @(posedge clk)
m0111111_1<=h0111111_1;
always @(posedge clk)
m1000000_0<=h1000000_0;
always @(posedge clk)
m1000000_1<=h1000000_1;
always @(posedge clk)
m1000001_0<=h1000001_0;
always @(posedge clk)
m1000001_1<=h1000001_1;
always @(posedge clk)
m1000010_0<=h1000010_0;
always @(posedge clk)
m1000010_1<=h1000010_1;
always @(posedge clk)
m1000011_0<=h1000011_0;
always @(posedge clk)
m1000011_1<=h1000011_1;
always @(posedge clk)
m1000100_0<=h1000100_0;
always @(posedge clk)
m1000100_1<=h1000100_1;
always @(posedge clk)
m1000101_0<=h1000101_0;
always @(posedge clk)
m1000101_1<=h1000101_1;
always @(posedge clk)
m1000110_0<=h1000110_0;
always @(posedge clk)
m1000110_1<=h1000110_1;
always @(posedge clk)
m1000111_0<=h1000111_0;
always @(posedge clk)
m1000111_1<=h1000111_1;
always @(posedge clk)
m1001000_0<=h1001000_0;
always @(posedge clk)
m1001000_1<=h1001000_1;
always @(posedge clk)
m1001001_0<=h1001001_0;
always @(posedge clk)
m1001001_1<=h1001001_1;
always @(posedge clk)
m1001010_0<=h1001010_0;
always @(posedge clk)
m1001010_1<=h1001010_1;
always @(posedge clk)
m1001011_0<=h1001011_0;
always @(posedge clk)
m1001011_1<=h1001011_1;
always @(posedge clk)
m1001100_0<=h1001100_0;
always @(posedge clk)
m1001100_1<=h1001100_1;
always @(posedge clk)
m1001101_0<=h1001101_0;
always @(posedge clk)
m1001101_1<=h1001101_1;
always @(posedge clk)
m1001110_0<=h1001110_0;
always @(posedge clk)
m1001110_1<=h1001110_1;
always @(posedge clk)
m1001111_0<=h1001111_0;
always @(posedge clk)
m1001111_1<=h1001111_1;
always @(posedge clk)
m1010000_0<=h1010000_0;
always @(posedge clk)
m1010000_1<=h1010000_1;
always @(posedge clk)
m1010001_0<=h1010001_0;
always @(posedge clk)
m1010001_1<=h1010001_1;
always @(posedge clk)
m1010010_0<=h1010010_0;
always @(posedge clk)
m1010010_1<=h1010010_1;
always @(posedge clk)
m1010011_0<=h1010011_0;
always @(posedge clk)
m1010011_1<=h1010011_1;
always @(posedge clk)
m1010100_0<=h1010100_0;
always @(posedge clk)
m1010100_1<=h1010100_1;
always @(posedge clk)
m1010101_0<=h1010101_0;
always @(posedge clk)
m1010101_1<=h1010101_1;
always @(posedge clk)
m1010110_0<=h1010110_0;
always @(posedge clk)
m1010110_1<=h1010110_1;
always @(posedge clk)
m1010111_0<=h1010111_0;
always @(posedge clk)
m1010111_1<=h1010111_1;
always @(posedge clk)
m1011000_0<=h1011000_0;
always @(posedge clk)
m1011000_1<=h1011000_1;
always @(posedge clk)
m1011001_0<=h1011001_0;
always @(posedge clk)
m1011001_1<=h1011001_1;
always @(posedge clk)
m1011010_0<=h1011010_0;
always @(posedge clk)
m1011010_1<=h1011010_1;
always @(posedge clk)
m1011011_0<=h1011011_0;
always @(posedge clk)
m1011011_1<=h1011011_1;
always @(posedge clk)
m1011100_0<=h1011100_0;
always @(posedge clk)
m1011100_1<=h1011100_1;
always @(posedge clk)
m1011101_0<=h1011101_0;
always @(posedge clk)
m1011101_1<=h1011101_1;
always @(posedge clk)
m1011110_0<=h1011110_0;
always @(posedge clk)
m1011110_1<=h1011110_1;
always @(posedge clk)
m1011111_0<=h1011111_0;
always @(posedge clk)
m1011111_1<=h1011111_1;
always @(posedge clk)
m1100000_0<=h1100000_0;
always @(posedge clk)
m1100000_1<=h1100000_1;
always @(posedge clk)
m1100001_0<=h1100001_0;
always @(posedge clk)
m1100001_1<=h1100001_1;
always @(posedge clk)
m1100010_0<=h1100010_0;
always @(posedge clk)
m1100010_1<=h1100010_1;
always @(posedge clk)
m1100011_0<=h1100011_0;
always @(posedge clk)
m1100011_1<=h1100011_1;
always @(posedge clk)
m1100100_0<=h1100100_0;
always @(posedge clk)
m1100100_1<=h1100100_1;
always @(posedge clk)
m1100101_0<=h1100101_0;
always @(posedge clk)
m1100101_1<=h1100101_1;
always @(posedge clk)
m1100110_0<=h1100110_0;
always @(posedge clk)
m1100110_1<=h1100110_1;
always @(posedge clk)
m1100111_0<=h1100111_0;
always @(posedge clk)
m1100111_1<=h1100111_1;
always @(posedge clk)
m1101000_0<=h1101000_0;
always @(posedge clk)
m1101000_1<=h1101000_1;
always @(posedge clk)
m1101001_0<=h1101001_0;
always @(posedge clk)
m1101001_1<=h1101001_1;
always @(posedge clk)
m1101010_0<=h1101010_0;
always @(posedge clk)
m1101010_1<=h1101010_1;
always @(posedge clk)
m1101011_0<=h1101011_0;
always @(posedge clk)
m1101011_1<=h1101011_1;
always @(posedge clk)
m1101100_0<=h1101100_0;
always @(posedge clk)
m1101100_1<=h1101100_1;
always @(posedge clk)
m1101101_0<=h1101101_0;
always @(posedge clk)
m1101101_1<=h1101101_1;
always @(posedge clk)
m1101110_0<=h1101110_0;
always @(posedge clk)
m1101110_1<=h1101110_1;
always @(posedge clk)
m1101111_0<=h1101111_0;
always @(posedge clk)
m1101111_1<=h1101111_1;
always @(posedge clk)
m1110000_0<=h1110000_0;
always @(posedge clk)
m1110000_1<=h1110000_1;
always @(posedge clk)
m1110001_0<=h1110001_0;
always @(posedge clk)
m1110001_1<=h1110001_1;
always @(posedge clk)
m1110010_0<=h1110010_0;
always @(posedge clk)
m1110010_1<=h1110010_1;
always @(posedge clk)
m1110011_0<=h1110011_0;
always @(posedge clk)
m1110011_1<=h1110011_1;
always @(posedge clk)
m1110100_0<=h1110100_0;
always @(posedge clk)
m1110100_1<=h1110100_1;
always @(posedge clk)
m1110101_0<=h1110101_0;
always @(posedge clk)
m1110101_1<=h1110101_1;
always @(posedge clk)
m1110110_0<=h1110110_0;
always @(posedge clk)
m1110110_1<=h1110110_1;
always @(posedge clk)
m1110111_0<=h1110111_0;
always @(posedge clk)
m1110111_1<=h1110111_1;
always @(posedge clk)
m1111000_0<=h1111000_0;
always @(posedge clk)
m1111000_1<=h1111000_1;
always @(posedge clk)
m1111001_0<=h1111001_0;
always @(posedge clk)
m1111001_1<=h1111001_1;
always @(posedge clk)
m1111010_0<=h1111010_0;
always @(posedge clk)
m1111010_1<=h1111010_1;
always @(posedge clk)
m1111011_0<=h1111011_0;
always @(posedge clk)
m1111011_1<=h1111011_1;
always @(posedge clk)
m1111100_0<=h1111100_0;
always @(posedge clk)
m1111100_1<=h1111100_1;
always @(posedge clk)
m1111101_0<=h1111101_0;
always @(posedge clk)
m1111101_1<=h1111101_1;
always @(posedge clk)
m1111110_0<=h1111110_0;
always @(posedge clk)
m1111110_1<=h1111110_1;
always @(posedge clk)
m1111111_0<=h1111111_0;
always @(posedge clk)
m1111111_1<=h1111111_1;

always @(negedge clk)
q0000000_0<=m0000000_0;
always @(negedge clk)
q0000000_1<=m0000000_1;
always @(negedge clk)
q0000001_0<=m0000001_0;
always @(negedge clk)
q0000001_1<=m0000001_1;
always @(negedge clk)
q0000010_0<=m0000010_0;
always @(negedge clk)
q0000010_1<=m0000010_1;
always @(negedge clk)
q0000011_0<=m0000011_0;
always @(negedge clk)
q0000011_1<=m0000011_1;
always @(negedge clk)
q0000100_0<=m0000100_0;
always @(negedge clk)
q0000100_1<=m0000100_1;
always @(negedge clk)
q0000101_0<=m0000101_0;
always @(negedge clk)
q0000101_1<=m0000101_1;
always @(negedge clk)
q0000110_0<=m0000110_0;
always @(negedge clk)
q0000110_1<=m0000110_1;
always @(negedge clk)
q0000111_0<=m0000111_0;
always @(negedge clk)
q0000111_1<=m0000111_1;
always @(negedge clk)
q0001000_0<=m0001000_0;
always @(negedge clk)
q0001000_1<=m0001000_1;
always @(negedge clk)
q0001001_0<=m0001001_0;
always @(negedge clk)
q0001001_1<=m0001001_1;
always @(negedge clk)
q0001010_0<=m0001010_0;
always @(negedge clk)
q0001010_1<=m0001010_1;
always @(negedge clk)
q0001011_0<=m0001011_0;
always @(negedge clk)
q0001011_1<=m0001011_1;
always @(negedge clk)
q0001100_0<=m0001100_0;
always @(negedge clk)
q0001100_1<=m0001100_1;
always @(negedge clk)
q0001101_0<=m0001101_0;
always @(negedge clk)
q0001101_1<=m0001101_1;
always @(negedge clk)
q0001110_0<=m0001110_0;
always @(negedge clk)
q0001110_1<=m0001110_1;
always @(negedge clk)
q0001111_0<=m0001111_0;
always @(negedge clk)
q0001111_1<=m0001111_1;
always @(negedge clk)
q0010000_0<=m0010000_0;
always @(negedge clk)
q0010000_1<=m0010000_1;
always @(negedge clk)
q0010001_0<=m0010001_0;
always @(negedge clk)
q0010001_1<=m0010001_1;
always @(negedge clk)
q0010010_0<=m0010010_0;
always @(negedge clk)
q0010010_1<=m0010010_1;
always @(negedge clk)
q0010011_0<=m0010011_0;
always @(negedge clk)
q0010011_1<=m0010011_1;
always @(negedge clk)
q0010100_0<=m0010100_0;
always @(negedge clk)
q0010100_1<=m0010100_1;
always @(negedge clk)
q0010101_0<=m0010101_0;
always @(negedge clk)
q0010101_1<=m0010101_1;
always @(negedge clk)
q0010110_0<=m0010110_0;
always @(negedge clk)
q0010110_1<=m0010110_1;
always @(negedge clk)
q0010111_0<=m0010111_0;
always @(negedge clk)
q0010111_1<=m0010111_1;
always @(negedge clk)
q0011000_0<=m0011000_0;
always @(negedge clk)
q0011000_1<=m0011000_1;
always @(negedge clk)
q0011001_0<=m0011001_0;
always @(negedge clk)
q0011001_1<=m0011001_1;
always @(negedge clk)
q0011010_0<=m0011010_0;
always @(negedge clk)
q0011010_1<=m0011010_1;
always @(negedge clk)
q0011011_0<=m0011011_0;
always @(negedge clk)
q0011011_1<=m0011011_1;
always @(negedge clk)
q0011100_0<=m0011100_0;
always @(negedge clk)
q0011100_1<=m0011100_1;
always @(negedge clk)
q0011101_0<=m0011101_0;
always @(negedge clk)
q0011101_1<=m0011101_1;
always @(negedge clk)
q0011110_0<=m0011110_0;
always @(negedge clk)
q0011110_1<=m0011110_1;
always @(negedge clk)
q0011111_0<=m0011111_0;
always @(negedge clk)
q0011111_1<=m0011111_1;
always @(negedge clk)
q0100000_0<=m0100000_0;
always @(negedge clk)
q0100000_1<=m0100000_1;
always @(negedge clk)
q0100001_0<=m0100001_0;
always @(negedge clk)
q0100001_1<=m0100001_1;
always @(negedge clk)
q0100010_0<=m0100010_0;
always @(negedge clk)
q0100010_1<=m0100010_1;
always @(negedge clk)
q0100011_0<=m0100011_0;
always @(negedge clk)
q0100011_1<=m0100011_1;
always @(negedge clk)
q0100100_0<=m0100100_0;
always @(negedge clk)
q0100100_1<=m0100100_1;
always @(negedge clk)
q0100101_0<=m0100101_0;
always @(negedge clk)
q0100101_1<=m0100101_1;
always @(negedge clk)
q0100110_0<=m0100110_0;
always @(negedge clk)
q0100110_1<=m0100110_1;
always @(negedge clk)
q0100111_0<=m0100111_0;
always @(negedge clk)
q0100111_1<=m0100111_1;
always @(negedge clk)
q0101000_0<=m0101000_0;
always @(negedge clk)
q0101000_1<=m0101000_1;
always @(negedge clk)
q0101001_0<=m0101001_0;
always @(negedge clk)
q0101001_1<=m0101001_1;
always @(negedge clk)
q0101010_0<=m0101010_0;
always @(negedge clk)
q0101010_1<=m0101010_1;
always @(negedge clk)
q0101011_0<=m0101011_0;
always @(negedge clk)
q0101011_1<=m0101011_1;
always @(negedge clk)
q0101100_0<=m0101100_0;
always @(negedge clk)
q0101100_1<=m0101100_1;
always @(negedge clk)
q0101101_0<=m0101101_0;
always @(negedge clk)
q0101101_1<=m0101101_1;
always @(negedge clk)
q0101110_0<=m0101110_0;
always @(negedge clk)
q0101110_1<=m0101110_1;
always @(negedge clk)
q0101111_0<=m0101111_0;
always @(negedge clk)
q0101111_1<=m0101111_1;
always @(negedge clk)
q0110000_0<=m0110000_0;
always @(negedge clk)
q0110000_1<=m0110000_1;
always @(negedge clk)
q0110001_0<=m0110001_0;
always @(negedge clk)
q0110001_1<=m0110001_1;
always @(negedge clk)
q0110010_0<=m0110010_0;
always @(negedge clk)
q0110010_1<=m0110010_1;
always @(negedge clk)
q0110011_0<=m0110011_0;
always @(negedge clk)
q0110011_1<=m0110011_1;
always @(negedge clk)
q0110100_0<=m0110100_0;
always @(negedge clk)
q0110100_1<=m0110100_1;
always @(negedge clk)
q0110101_0<=m0110101_0;
always @(negedge clk)
q0110101_1<=m0110101_1;
always @(negedge clk)
q0110110_0<=m0110110_0;
always @(negedge clk)
q0110110_1<=m0110110_1;
always @(negedge clk)
q0110111_0<=m0110111_0;
always @(negedge clk)
q0110111_1<=m0110111_1;
always @(negedge clk)
q0111000_0<=m0111000_0;
always @(negedge clk)
q0111000_1<=m0111000_1;
always @(negedge clk)
q0111001_0<=m0111001_0;
always @(negedge clk)
q0111001_1<=m0111001_1;
always @(negedge clk)
q0111010_0<=m0111010_0;
always @(negedge clk)
q0111010_1<=m0111010_1;
always @(negedge clk)
q0111011_0<=m0111011_0;
always @(negedge clk)
q0111011_1<=m0111011_1;
always @(negedge clk)
q0111100_0<=m0111100_0;
always @(negedge clk)
q0111100_1<=m0111100_1;
always @(negedge clk)
q0111101_0<=m0111101_0;
always @(negedge clk)
q0111101_1<=m0111101_1;
always @(negedge clk)
q0111110_0<=m0111110_0;
always @(negedge clk)
q0111110_1<=m0111110_1;
always @(negedge clk)
q0111111_0<=m0111111_0;
always @(negedge clk)
q0111111_1<=m0111111_1;
always @(negedge clk)
q1000000_0<=m1000000_0;
always @(negedge clk)
q1000000_1<=m1000000_1;
always @(negedge clk)
q1000001_0<=m1000001_0;
always @(negedge clk)
q1000001_1<=m1000001_1;
always @(negedge clk)
q1000010_0<=m1000010_0;
always @(negedge clk)
q1000010_1<=m1000010_1;
always @(negedge clk)
q1000011_0<=m1000011_0;
always @(negedge clk)
q1000011_1<=m1000011_1;
always @(negedge clk)
q1000100_0<=m1000100_0;
always @(negedge clk)
q1000100_1<=m1000100_1;
always @(negedge clk)
q1000101_0<=m1000101_0;
always @(negedge clk)
q1000101_1<=m1000101_1;
always @(negedge clk)
q1000110_0<=m1000110_0;
always @(negedge clk)
q1000110_1<=m1000110_1;
always @(negedge clk)
q1000111_0<=m1000111_0;
always @(negedge clk)
q1000111_1<=m1000111_1;
always @(negedge clk)
q1001000_0<=m1001000_0;
always @(negedge clk)
q1001000_1<=m1001000_1;
always @(negedge clk)
q1001001_0<=m1001001_0;
always @(negedge clk)
q1001001_1<=m1001001_1;
always @(negedge clk)
q1001010_0<=m1001010_0;
always @(negedge clk)
q1001010_1<=m1001010_1;
always @(negedge clk)
q1001011_0<=m1001011_0;
always @(negedge clk)
q1001011_1<=m1001011_1;
always @(negedge clk)
q1001100_0<=m1001100_0;
always @(negedge clk)
q1001100_1<=m1001100_1;
always @(negedge clk)
q1001101_0<=m1001101_0;
always @(negedge clk)
q1001101_1<=m1001101_1;
always @(negedge clk)
q1001110_0<=m1001110_0;
always @(negedge clk)
q1001110_1<=m1001110_1;
always @(negedge clk)
q1001111_0<=m1001111_0;
always @(negedge clk)
q1001111_1<=m1001111_1;
always @(negedge clk)
q1010000_0<=m1010000_0;
always @(negedge clk)
q1010000_1<=m1010000_1;
always @(negedge clk)
q1010001_0<=m1010001_0;
always @(negedge clk)
q1010001_1<=m1010001_1;
always @(negedge clk)
q1010010_0<=m1010010_0;
always @(negedge clk)
q1010010_1<=m1010010_1;
always @(negedge clk)
q1010011_0<=m1010011_0;
always @(negedge clk)
q1010011_1<=m1010011_1;
always @(negedge clk)
q1010100_0<=m1010100_0;
always @(negedge clk)
q1010100_1<=m1010100_1;
always @(negedge clk)
q1010101_0<=m1010101_0;
always @(negedge clk)
q1010101_1<=m1010101_1;
always @(negedge clk)
q1010110_0<=m1010110_0;
always @(negedge clk)
q1010110_1<=m1010110_1;
always @(negedge clk)
q1010111_0<=m1010111_0;
always @(negedge clk)
q1010111_1<=m1010111_1;
always @(negedge clk)
q1011000_0<=m1011000_0;
always @(negedge clk)
q1011000_1<=m1011000_1;
always @(negedge clk)
q1011001_0<=m1011001_0;
always @(negedge clk)
q1011001_1<=m1011001_1;
always @(negedge clk)
q1011010_0<=m1011010_0;
always @(negedge clk)
q1011010_1<=m1011010_1;
always @(negedge clk)
q1011011_0<=m1011011_0;
always @(negedge clk)
q1011011_1<=m1011011_1;
always @(negedge clk)
q1011100_0<=m1011100_0;
always @(negedge clk)
q1011100_1<=m1011100_1;
always @(negedge clk)
q1011101_0<=m1011101_0;
always @(negedge clk)
q1011101_1<=m1011101_1;
always @(negedge clk)
q1011110_0<=m1011110_0;
always @(negedge clk)
q1011110_1<=m1011110_1;
always @(negedge clk)
q1011111_0<=m1011111_0;
always @(negedge clk)
q1011111_1<=m1011111_1;
always @(negedge clk)
q1100000_0<=m1100000_0;
always @(negedge clk)
q1100000_1<=m1100000_1;
always @(negedge clk)
q1100001_0<=m1100001_0;
always @(negedge clk)
q1100001_1<=m1100001_1;
always @(negedge clk)
q1100010_0<=m1100010_0;
always @(negedge clk)
q1100010_1<=m1100010_1;
always @(negedge clk)
q1100011_0<=m1100011_0;
always @(negedge clk)
q1100011_1<=m1100011_1;
always @(negedge clk)
q1100100_0<=m1100100_0;
always @(negedge clk)
q1100100_1<=m1100100_1;
always @(negedge clk)
q1100101_0<=m1100101_0;
always @(negedge clk)
q1100101_1<=m1100101_1;
always @(negedge clk)
q1100110_0<=m1100110_0;
always @(negedge clk)
q1100110_1<=m1100110_1;
always @(negedge clk)
q1100111_0<=m1100111_0;
always @(negedge clk)
q1100111_1<=m1100111_1;
always @(negedge clk)
q1101000_0<=m1101000_0;
always @(negedge clk)
q1101000_1<=m1101000_1;
always @(negedge clk)
q1101001_0<=m1101001_0;
always @(negedge clk)
q1101001_1<=m1101001_1;
always @(negedge clk)
q1101010_0<=m1101010_0;
always @(negedge clk)
q1101010_1<=m1101010_1;
always @(negedge clk)
q1101011_0<=m1101011_0;
always @(negedge clk)
q1101011_1<=m1101011_1;
always @(negedge clk)
q1101100_0<=m1101100_0;
always @(negedge clk)
q1101100_1<=m1101100_1;
always @(negedge clk)
q1101101_0<=m1101101_0;
always @(negedge clk)
q1101101_1<=m1101101_1;
always @(negedge clk)
q1101110_0<=m1101110_0;
always @(negedge clk)
q1101110_1<=m1101110_1;
always @(negedge clk)
q1101111_0<=m1101111_0;
always @(negedge clk)
q1101111_1<=m1101111_1;
always @(negedge clk)
q1110000_0<=m1110000_0;
always @(negedge clk)
q1110000_1<=m1110000_1;
always @(negedge clk)
q1110001_0<=m1110001_0;
always @(negedge clk)
q1110001_1<=m1110001_1;
always @(negedge clk)
q1110010_0<=m1110010_0;
always @(negedge clk)
q1110010_1<=m1110010_1;
always @(negedge clk)
q1110011_0<=m1110011_0;
always @(negedge clk)
q1110011_1<=m1110011_1;
always @(negedge clk)
q1110100_0<=m1110100_0;
always @(negedge clk)
q1110100_1<=m1110100_1;
always @(negedge clk)
q1110101_0<=m1110101_0;
always @(negedge clk)
q1110101_1<=m1110101_1;
always @(negedge clk)
q1110110_0<=m1110110_0;
always @(negedge clk)
q1110110_1<=m1110110_1;
always @(negedge clk)
q1110111_0<=m1110111_0;
always @(negedge clk)
q1110111_1<=m1110111_1;
always @(negedge clk)
q1111000_0<=m1111000_0;
always @(negedge clk)
q1111000_1<=m1111000_1;
always @(negedge clk)
q1111001_0<=m1111001_0;
always @(negedge clk)
q1111001_1<=m1111001_1;
always @(negedge clk)
q1111010_0<=m1111010_0;
always @(negedge clk)
q1111010_1<=m1111010_1;
always @(negedge clk)
q1111011_0<=m1111011_0;
always @(negedge clk)
q1111011_1<=m1111011_1;
always @(negedge clk)
q1111100_0<=m1111100_0;
always @(negedge clk)
q1111100_1<=m1111100_1;
always @(negedge clk)
q1111101_0<=m1111101_0;
always @(negedge clk)
q1111101_1<=m1111101_1;
always @(negedge clk)
q1111110_0<=m1111110_0;
always @(negedge clk)
q1111110_1<=m1111110_1;
always @(negedge clk)
q1111111_0<=m1111111_0;
always @(negedge clk)
q1111111_1<=m1111111_1;

always @(posedge clk)
m000000_0<=h000000_0;
always @(posedge clk)
m000000_1<=h000000_1;
always @(posedge clk)
m000001_0<=h000001_0;
always @(posedge clk)
m000001_1<=h000001_1;
always @(posedge clk)
m000010_0<=h000010_0;
always @(posedge clk)
m000010_1<=h000010_1;
always @(posedge clk)
m000011_0<=h000011_0;
always @(posedge clk)
m000011_1<=h000011_1;
always @(posedge clk)
m000100_0<=h000100_0;
always @(posedge clk)
m000100_1<=h000100_1;
always @(posedge clk)
m000101_0<=h000101_0;
always @(posedge clk)
m000101_1<=h000101_1;
always @(posedge clk)
m000110_0<=h000110_0;
always @(posedge clk)
m000110_1<=h000110_1;
always @(posedge clk)
m000111_0<=h000111_0;
always @(posedge clk)
m000111_1<=h000111_1;
always @(posedge clk)
m001000_0<=h001000_0;
always @(posedge clk)
m001000_1<=h001000_1;
always @(posedge clk)
m001001_0<=h001001_0;
always @(posedge clk)
m001001_1<=h001001_1;
always @(posedge clk)
m001010_0<=h001010_0;
always @(posedge clk)
m001010_1<=h001010_1;
always @(posedge clk)
m001011_0<=h001011_0;
always @(posedge clk)
m001011_1<=h001011_1;
always @(posedge clk)
m001100_0<=h001100_0;
always @(posedge clk)
m001100_1<=h001100_1;
always @(posedge clk)
m001101_0<=h001101_0;
always @(posedge clk)
m001101_1<=h001101_1;
always @(posedge clk)
m001110_0<=h001110_0;
always @(posedge clk)
m001110_1<=h001110_1;
always @(posedge clk)
m001111_0<=h001111_0;
always @(posedge clk)
m001111_1<=h001111_1;
always @(posedge clk)
m010000_0<=h010000_0;
always @(posedge clk)
m010000_1<=h010000_1;
always @(posedge clk)
m010001_0<=h010001_0;
always @(posedge clk)
m010001_1<=h010001_1;
always @(posedge clk)
m010010_0<=h010010_0;
always @(posedge clk)
m010010_1<=h010010_1;
always @(posedge clk)
m010011_0<=h010011_0;
always @(posedge clk)
m010011_1<=h010011_1;
always @(posedge clk)
m010100_0<=h010100_0;
always @(posedge clk)
m010100_1<=h010100_1;
always @(posedge clk)
m010101_0<=h010101_0;
always @(posedge clk)
m010101_1<=h010101_1;
always @(posedge clk)
m010110_0<=h010110_0;
always @(posedge clk)
m010110_1<=h010110_1;
always @(posedge clk)
m010111_0<=h010111_0;
always @(posedge clk)
m010111_1<=h010111_1;
always @(posedge clk)
m011000_0<=h011000_0;
always @(posedge clk)
m011000_1<=h011000_1;
always @(posedge clk)
m011001_0<=h011001_0;
always @(posedge clk)
m011001_1<=h011001_1;
always @(posedge clk)
m011010_0<=h011010_0;
always @(posedge clk)
m011010_1<=h011010_1;
always @(posedge clk)
m011011_0<=h011011_0;
always @(posedge clk)
m011011_1<=h011011_1;
always @(posedge clk)
m011100_0<=h011100_0;
always @(posedge clk)
m011100_1<=h011100_1;
always @(posedge clk)
m011101_0<=h011101_0;
always @(posedge clk)
m011101_1<=h011101_1;
always @(posedge clk)
m011110_0<=h011110_0;
always @(posedge clk)
m011110_1<=h011110_1;
always @(posedge clk)
m011111_0<=h011111_0;
always @(posedge clk)
m011111_1<=h011111_1;
always @(posedge clk)
m100000_0<=h100000_0;
always @(posedge clk)
m100000_1<=h100000_1;
always @(posedge clk)
m100001_0<=h100001_0;
always @(posedge clk)
m100001_1<=h100001_1;
always @(posedge clk)
m100010_0<=h100010_0;
always @(posedge clk)
m100010_1<=h100010_1;
always @(posedge clk)
m100011_0<=h100011_0;
always @(posedge clk)
m100011_1<=h100011_1;
always @(posedge clk)
m100100_0<=h100100_0;
always @(posedge clk)
m100100_1<=h100100_1;
always @(posedge clk)
m100101_0<=h100101_0;
always @(posedge clk)
m100101_1<=h100101_1;
always @(posedge clk)
m100110_0<=h100110_0;
always @(posedge clk)
m100110_1<=h100110_1;
always @(posedge clk)
m100111_0<=h100111_0;
always @(posedge clk)
m100111_1<=h100111_1;
always @(posedge clk)
m101000_0<=h101000_0;
always @(posedge clk)
m101000_1<=h101000_1;
always @(posedge clk)
m101001_0<=h101001_0;
always @(posedge clk)
m101001_1<=h101001_1;
always @(posedge clk)
m101010_0<=h101010_0;
always @(posedge clk)
m101010_1<=h101010_1;
always @(posedge clk)
m101011_0<=h101011_0;
always @(posedge clk)
m101011_1<=h101011_1;
always @(posedge clk)
m101100_0<=h101100_0;
always @(posedge clk)
m101100_1<=h101100_1;
always @(posedge clk)
m101101_0<=h101101_0;
always @(posedge clk)
m101101_1<=h101101_1;
always @(posedge clk)
m101110_0<=h101110_0;
always @(posedge clk)
m101110_1<=h101110_1;
always @(posedge clk)
m101111_0<=h101111_0;
always @(posedge clk)
m101111_1<=h101111_1;
always @(posedge clk)
m110000_0<=h110000_0;
always @(posedge clk)
m110000_1<=h110000_1;
always @(posedge clk)
m110001_0<=h110001_0;
always @(posedge clk)
m110001_1<=h110001_1;
always @(posedge clk)
m110010_0<=h110010_0;
always @(posedge clk)
m110010_1<=h110010_1;
always @(posedge clk)
m110011_0<=h110011_0;
always @(posedge clk)
m110011_1<=h110011_1;
always @(posedge clk)
m110100_0<=h110100_0;
always @(posedge clk)
m110100_1<=h110100_1;
always @(posedge clk)
m110101_0<=h110101_0;
always @(posedge clk)
m110101_1<=h110101_1;
always @(posedge clk)
m110110_0<=h110110_0;
always @(posedge clk)
m110110_1<=h110110_1;
always @(posedge clk)
m110111_0<=h110111_0;
always @(posedge clk)
m110111_1<=h110111_1;
always @(posedge clk)
m111000_0<=h111000_0;
always @(posedge clk)
m111000_1<=h111000_1;
always @(posedge clk)
m111001_0<=h111001_0;
always @(posedge clk)
m111001_1<=h111001_1;
always @(posedge clk)
m111010_0<=h111010_0;
always @(posedge clk)
m111010_1<=h111010_1;
always @(posedge clk)
m111011_0<=h111011_0;
always @(posedge clk)
m111011_1<=h111011_1;
always @(posedge clk)
m111100_0<=h111100_0;
always @(posedge clk)
m111100_1<=h111100_1;
always @(posedge clk)
m111101_0<=h111101_0;
always @(posedge clk)
m111101_1<=h111101_1;
always @(posedge clk)
m111110_0<=h111110_0;
always @(posedge clk)
m111110_1<=h111110_1;
always @(posedge clk)
m111111_0<=h111111_0;
always @(posedge clk)
m111111_1<=h111111_1;

always @(negedge clk)
q000000_0<=m000000_0;
always @(negedge clk)
q000000_1<=m000000_1;
always @(negedge clk)
q000001_0<=m000001_0;
always @(negedge clk)
q000001_1<=m000001_1;
always @(negedge clk)
q000010_0<=m000010_0;
always @(negedge clk)
q000010_1<=m000010_1;
always @(negedge clk)
q000011_0<=m000011_0;
always @(negedge clk)
q000011_1<=m000011_1;
always @(negedge clk)
q000100_0<=m000100_0;
always @(negedge clk)
q000100_1<=m000100_1;
always @(negedge clk)
q000101_0<=m000101_0;
always @(negedge clk)
q000101_1<=m000101_1;
always @(negedge clk)
q000110_0<=m000110_0;
always @(negedge clk)
q000110_1<=m000110_1;
always @(negedge clk)
q000111_0<=m000111_0;
always @(negedge clk)
q000111_1<=m000111_1;
always @(negedge clk)
q001000_0<=m001000_0;
always @(negedge clk)
q001000_1<=m001000_1;
always @(negedge clk)
q001001_0<=m001001_0;
always @(negedge clk)
q001001_1<=m001001_1;
always @(negedge clk)
q001010_0<=m001010_0;
always @(negedge clk)
q001010_1<=m001010_1;
always @(negedge clk)
q001011_0<=m001011_0;
always @(negedge clk)
q001011_1<=m001011_1;
always @(negedge clk)
q001100_0<=m001100_0;
always @(negedge clk)
q001100_1<=m001100_1;
always @(negedge clk)
q001101_0<=m001101_0;
always @(negedge clk)
q001101_1<=m001101_1;
always @(negedge clk)
q001110_0<=m001110_0;
always @(negedge clk)
q001110_1<=m001110_1;
always @(negedge clk)
q001111_0<=m001111_0;
always @(negedge clk)
q001111_1<=m001111_1;
always @(negedge clk)
q010000_0<=m010000_0;
always @(negedge clk)
q010000_1<=m010000_1;
always @(negedge clk)
q010001_0<=m010001_0;
always @(negedge clk)
q010001_1<=m010001_1;
always @(negedge clk)
q010010_0<=m010010_0;
always @(negedge clk)
q010010_1<=m010010_1;
always @(negedge clk)
q010011_0<=m010011_0;
always @(negedge clk)
q010011_1<=m010011_1;
always @(negedge clk)
q010100_0<=m010100_0;
always @(negedge clk)
q010100_1<=m010100_1;
always @(negedge clk)
q010101_0<=m010101_0;
always @(negedge clk)
q010101_1<=m010101_1;
always @(negedge clk)
q010110_0<=m010110_0;
always @(negedge clk)
q010110_1<=m010110_1;
always @(negedge clk)
q010111_0<=m010111_0;
always @(negedge clk)
q010111_1<=m010111_1;
always @(negedge clk)
q011000_0<=m011000_0;
always @(negedge clk)
q011000_1<=m011000_1;
always @(negedge clk)
q011001_0<=m011001_0;
always @(negedge clk)
q011001_1<=m011001_1;
always @(negedge clk)
q011010_0<=m011010_0;
always @(negedge clk)
q011010_1<=m011010_1;
always @(negedge clk)
q011011_0<=m011011_0;
always @(negedge clk)
q011011_1<=m011011_1;
always @(negedge clk)
q011100_0<=m011100_0;
always @(negedge clk)
q011100_1<=m011100_1;
always @(negedge clk)
q011101_0<=m011101_0;
always @(negedge clk)
q011101_1<=m011101_1;
always @(negedge clk)
q011110_0<=m011110_0;
always @(negedge clk)
q011110_1<=m011110_1;
always @(negedge clk)
q011111_0<=m011111_0;
always @(negedge clk)
q011111_1<=m011111_1;
always @(negedge clk)
q100000_0<=m100000_0;
always @(negedge clk)
q100000_1<=m100000_1;
always @(negedge clk)
q100001_0<=m100001_0;
always @(negedge clk)
q100001_1<=m100001_1;
always @(negedge clk)
q100010_0<=m100010_0;
always @(negedge clk)
q100010_1<=m100010_1;
always @(negedge clk)
q100011_0<=m100011_0;
always @(negedge clk)
q100011_1<=m100011_1;
always @(negedge clk)
q100100_0<=m100100_0;
always @(negedge clk)
q100100_1<=m100100_1;
always @(negedge clk)
q100101_0<=m100101_0;
always @(negedge clk)
q100101_1<=m100101_1;
always @(negedge clk)
q100110_0<=m100110_0;
always @(negedge clk)
q100110_1<=m100110_1;
always @(negedge clk)
q100111_0<=m100111_0;
always @(negedge clk)
q100111_1<=m100111_1;
always @(negedge clk)
q101000_0<=m101000_0;
always @(negedge clk)
q101000_1<=m101000_1;
always @(negedge clk)
q101001_0<=m101001_0;
always @(negedge clk)
q101001_1<=m101001_1;
always @(negedge clk)
q101010_0<=m101010_0;
always @(negedge clk)
q101010_1<=m101010_1;
always @(negedge clk)
q101011_0<=m101011_0;
always @(negedge clk)
q101011_1<=m101011_1;
always @(negedge clk)
q101100_0<=m101100_0;
always @(negedge clk)
q101100_1<=m101100_1;
always @(negedge clk)
q101101_0<=m101101_0;
always @(negedge clk)
q101101_1<=m101101_1;
always @(negedge clk)
q101110_0<=m101110_0;
always @(negedge clk)
q101110_1<=m101110_1;
always @(negedge clk)
q101111_0<=m101111_0;
always @(negedge clk)
q101111_1<=m101111_1;
always @(negedge clk)
q110000_0<=m110000_0;
always @(negedge clk)
q110000_1<=m110000_1;
always @(negedge clk)
q110001_0<=m110001_0;
always @(negedge clk)
q110001_1<=m110001_1;
always @(negedge clk)
q110010_0<=m110010_0;
always @(negedge clk)
q110010_1<=m110010_1;
always @(negedge clk)
q110011_0<=m110011_0;
always @(negedge clk)
q110011_1<=m110011_1;
always @(negedge clk)
q110100_0<=m110100_0;
always @(negedge clk)
q110100_1<=m110100_1;
always @(negedge clk)
q110101_0<=m110101_0;
always @(negedge clk)
q110101_1<=m110101_1;
always @(negedge clk)
q110110_0<=m110110_0;
always @(negedge clk)
q110110_1<=m110110_1;
always @(negedge clk)
q110111_0<=m110111_0;
always @(negedge clk)
q110111_1<=m110111_1;
always @(negedge clk)
q111000_0<=m111000_0;
always @(negedge clk)
q111000_1<=m111000_1;
always @(negedge clk)
q111001_0<=m111001_0;
always @(negedge clk)
q111001_1<=m111001_1;
always @(negedge clk)
q111010_0<=m111010_0;
always @(negedge clk)
q111010_1<=m111010_1;
always @(negedge clk)
q111011_0<=m111011_0;
always @(negedge clk)
q111011_1<=m111011_1;
always @(negedge clk)
q111100_0<=m111100_0;
always @(negedge clk)
q111100_1<=m111100_1;
always @(negedge clk)
q111101_0<=m111101_0;
always @(negedge clk)
q111101_1<=m111101_1;
always @(negedge clk)
q111110_0<=m111110_0;
always @(negedge clk)
q111110_1<=m111110_1;
always @(negedge clk)
q111111_0<=m111111_0;
always @(negedge clk)
q111111_1<=m111111_1;

always @(posedge clk)
m0001<=n0001;
always @(posedge clk)
m0002<=x0002;
always @(posedge clk)
m0003<=x0003;
always @(posedge clk)
m0004<=x0004;
always @(posedge clk)
m0005<=x0005;
always @(posedge clk)
m0006<=x0006;
always @(posedge clk)
m0007<=x0007;
always @(posedge clk)
m0008<=x0008;
always @(posedge clk)
m0009<=x0009;
always @(posedge clk)
m0010<=x0010;
always @(posedge clk)
m0011<=x0011;
always @(posedge clk)
m0012<=x0012;
always @(posedge clk)
m0013<=x0013;
always @(posedge clk)
m0014<=x0014;
always @(posedge clk)
m0015<=x0015;
always @(posedge clk)
m0016<=x0016;
always @(posedge clk)
m0017<=x0017;
always @(posedge clk)
m0018<=x0018;
always @(posedge clk)
m0019<=x0019;
always @(posedge clk)
m0020<=x0020;
always @(posedge clk)
m0021<=x0021;
always @(posedge clk)
m0022<=x0022;
always @(posedge clk)
m0023<=x0023;
always @(posedge clk)
m0024<=x0024;
always @(posedge clk)
m0025<=x0025;
always @(posedge clk)
m0026<=x0026;
always @(posedge clk)
m0027<=x0027;
always @(posedge clk)
m0028<=x0028;
always @(posedge clk)
m0029<=x0029;
always @(posedge clk)
m0030<=x0030;

always @(negedge clk)
q0001<=m0001;
always @(negedge clk)
q0002<=m0002;
always @(negedge clk)
q0003<=m0003;
always @(negedge clk)
q0004<=m0004;
always @(negedge clk)
q0005<=m0005;
always @(negedge clk)
q0006<=m0006;
always @(negedge clk)
q0007<=m0007;
always @(negedge clk)
q0008<=m0008;
always @(negedge clk)
q0009<=m0009;
always @(negedge clk)
q0010<=m0010;
always @(negedge clk)
q0011<=m0011;
always @(negedge clk)
q0012<=m0012;
always @(negedge clk)
q0013<=m0013;
always @(negedge clk)
q0014<=m0014;
always @(negedge clk)
q0015<=m0015;
always @(negedge clk)
q0016<=m0016;
always @(negedge clk)
q0017<=m0017;
always @(negedge clk)
q0018<=m0018;
always @(negedge clk)
q0019<=m0019;
always @(negedge clk)
q0020<=m0020;
always @(negedge clk)
q0021<=m0021;
always @(negedge clk)
q0022<=m0022;
always @(negedge clk)
q0023<=m0023;
always @(negedge clk)
q0024<=m0024;
always @(negedge clk)
q0025<=m0025;
always @(negedge clk)
q0026<=m0026;
always @(negedge clk)
q0027<=m0027;
always @(negedge clk)
q0028<=m0028;
always @(negedge clk)
q0029<=m0029;
always @(negedge clk)
q0030<=m0030;
//x
always @(posedge clk)
m0031<=a0061;
always @(posedge clk)
m0032<=a0062;
always @(posedge clk)
m0033<=a0063;
always @(posedge clk)
m0034<=a0064;
always @(posedge clk)
m0035<=a0065;
always @(posedge clk)
m0036<=a0066;
always @(posedge clk)
m0037<=a0067;
always @(posedge clk)
m0038<=a0068;
always @(posedge clk)
m0039<=a0069;
always @(posedge clk)
m0040<=a0070;
always @(posedge clk)
m0041<=a0071;
always @(posedge clk)
m0042<=a0072;
always @(posedge clk)
m0043<=a0073;
always @(posedge clk)
m0044<=a0074;
always @(posedge clk)
m0045<=a0075;
always @(posedge clk)
m0046<=a0076;
always @(posedge clk)
m0047<=a0077;
always @(posedge clk)
m0048<=a0078;
always @(posedge clk)
m0049<=a0079;
always @(posedge clk)
m0050<=a0080;
always @(posedge clk)
m0051<=a0081;
always @(posedge clk)
m0052<=a0082;
always @(posedge clk)
m0053<=a0083;
always @(posedge clk)
m0054<=a0084;
always @(posedge clk)
m0055<=a0085;
always @(posedge clk)
m0056<=a0086;
always @(posedge clk)
m0057<=a0087;
always @(posedge clk)
m0058<=a0088;
always @(posedge clk)
m0059<=a0089;
always @(posedge clk)
m0060<=a0090;

always @(negedge clk)
q0031<=m0031;
always @(negedge clk)
q0032<=m0032;
always @(negedge clk)
q0033<=m0033;
always @(negedge clk)
q0034<=m0034;
always @(negedge clk)
q0035<=m0035;
always @(negedge clk)
q0036<=m0036;
always @(negedge clk)
q0037<=m0037;
always @(negedge clk)
q0038<=m0038;
always @(negedge clk)
q0039<=m0039;
always @(negedge clk)
q0040<=m0040;
always @(negedge clk)
q0041<=m0041;
always @(negedge clk)
q0042<=m0042;
always @(negedge clk)
q0043<=m0043;
always @(negedge clk)
q0044<=m0044;
always @(negedge clk)
q0045<=m0045;
always @(negedge clk)
q0046<=m0046;
always @(negedge clk)
q0047<=m0047;
always @(negedge clk)
q0048<=m0048;
always @(negedge clk)
q0049<=m0049;
always @(negedge clk)
q0050<=m0050;
always @(negedge clk)
q0051<=m0051;
always @(negedge clk)
q0052<=m0052;
always @(negedge clk)
q0053<=m0053;
always @(negedge clk)
q0054<=m0054;
always @(negedge clk)
q0055<=m0055;
always @(negedge clk)
q0056<=m0056;
always @(negedge clk)
q0057<=m0057;
always @(negedge clk)
q0058<=m0058;
always @(negedge clk)
q0059<=m0059;
always @(negedge clk)
q0060<=m0060;

always @(posedge clk)
m0061<=h006101;
always @(posedge clk)
m0062<=h006201;
always @(posedge clk)
m0063<=h006301;
always @(posedge clk)
m0064<=h006401;
always @(posedge clk)
m0065<=h006501;
always @(posedge clk)
m0066<=h006601;
always @(posedge clk)
m0067<=h006701;
always @(posedge clk)
m0068<=h006801;
always @(posedge clk)
m0069<=h006901;
always @(posedge clk)
m0070<=h007001;
always @(posedge clk)
m0071<=h007101;
always @(posedge clk)
m0072<=h007201;
always @(posedge clk)
m0073<=h007301;
always @(posedge clk)
m0074<=h007401;
always @(posedge clk)
m0075<=h007501;
always @(posedge clk)
m0076<=h007601;
always @(posedge clk)
m0077<=h007701;
always @(posedge clk)
m0078<=h007801;
always @(posedge clk)
m0079<=h007901;
always @(posedge clk)
m0080<=h008001;
always @(posedge clk)
m0081<=h008101;
always @(posedge clk)
m0082<=h008201;
always @(posedge clk)
m0083<=h008301;
always @(posedge clk)
m0084<=h008401;
always @(posedge clk)
m0085<=h008501;
always @(posedge clk)
m0086<=h008601;
always @(posedge clk)
m0087<=h008701;
always @(posedge clk)
m0088<=h008801;
always @(posedge clk)
m0089<=h008901;
always @(posedge clk)
m0090<=h009001;

always @(negedge clk)
q0061<=m0061;
always @(negedge clk)
q0062<=m0062;
always @(negedge clk)
q0063<=m0063;
always @(negedge clk)
q0064<=m0064;
always @(negedge clk)
q0065<=m0065;
always @(negedge clk)
q0066<=m0066;
always @(negedge clk)
q0067<=m0067;
always @(negedge clk)
q0068<=m0068;
always @(negedge clk)
q0069<=m0069;
always @(negedge clk)
q0070<=m0070;
always @(negedge clk)
q0071<=m0071;
always @(negedge clk)
q0072<=m0072;
always @(negedge clk)
q0073<=m0073;
always @(negedge clk)
q0074<=m0074;
always @(negedge clk)
q0075<=m0075;
always @(negedge clk)
q0076<=m0076;
always @(negedge clk)
q0077<=m0077;
always @(negedge clk)
q0078<=m0078;
always @(negedge clk)
q0079<=m0079;
always @(negedge clk)
q0080<=m0080;
always @(negedge clk)
q0081<=m0081;
always @(negedge clk)
q0082<=m0082;
always @(negedge clk)
q0083<=m0083;
always @(negedge clk)
q0084<=m0084;
always @(negedge clk)
q0085<=m0085;
always @(negedge clk)
q0086<=m0086;
always @(negedge clk)
q0087<=m0087;
always @(negedge clk)
q0088<=m0088;
always @(negedge clk)
q0089<=m0089;
always @(negedge clk)
q0090<=m0090;
//y
always @(posedge clk)
m0091<=a0121;
always @(posedge clk)
m0092<=a0122;
always @(posedge clk)
m0093<=a0123;
always @(posedge clk)
m0094<=a0124;
always @(posedge clk)
m0095<=a0125;
always @(posedge clk)
m0096<=a0126;
always @(posedge clk)
m0097<=a0127;
always @(posedge clk)
m0098<=a0128;
always @(posedge clk)
m0099<=a0129;
always @(posedge clk)
m0100<=a0130;
always @(posedge clk)
m0101<=a0131;
always @(posedge clk)
m0102<=a0132;
always @(posedge clk)
m0103<=a0133;
always @(posedge clk)
m0104<=a0134;
always @(posedge clk)
m0105<=a0135;
always @(posedge clk)
m0106<=a0136;
always @(posedge clk)
m0107<=a0137;
always @(posedge clk)
m0108<=a0138;
always @(posedge clk)
m0109<=a0139;
always @(posedge clk)
m0110<=a0140;
always @(posedge clk)
m0111<=a0141;
always @(posedge clk)
m0112<=a0142;
always @(posedge clk)
m0113<=a0143;
always @(posedge clk)
m0114<=a0144;
always @(posedge clk)
m0115<=a0145;
always @(posedge clk)
m0116<=a0146;
always @(posedge clk)
m0117<=a0147;
always @(posedge clk)
m0118<=a0148;
always @(posedge clk)
m0119<=a0149;
always @(posedge clk)
m0120<=a0150;

always @(negedge clk)
q0091<=m0091;
always @(negedge clk)
q0092<=m0092;
always @(negedge clk)
q0093<=m0093;
always @(negedge clk)
q0094<=m0094;
always @(negedge clk)
q0095<=m0095;
always @(negedge clk)
q0096<=m0096;
always @(negedge clk)
q0097<=m0097;
always @(negedge clk)
q0098<=m0098;
always @(negedge clk)
q0099<=m0099;
always @(negedge clk)
q0100<=m0100;
always @(negedge clk)
q0101<=m0101;
always @(negedge clk)
q0102<=m0102;
always @(negedge clk)
q0103<=m0103;
always @(negedge clk)
q0104<=m0104;
always @(negedge clk)
q0105<=m0105;
always @(negedge clk)
q0106<=m0106;
always @(negedge clk)
q0107<=m0107;
always @(negedge clk)
q0108<=m0108;
always @(negedge clk)
q0109<=m0109;
always @(negedge clk)
q0110<=m0110;
always @(negedge clk)
q0111<=m0111;
always @(negedge clk)
q0112<=m0112;
always @(negedge clk)
q0113<=m0113;
always @(negedge clk)
q0114<=m0114;
always @(negedge clk)
q0115<=m0115;
always @(negedge clk)
q0116<=m0116;
always @(negedge clk)
q0117<=m0117;
always @(negedge clk)
q0118<=m0118;
always @(negedge clk)
q0119<=m0119;
always @(negedge clk)
q0120<=m0120;

always @(posedge clk)
m0121<=h012101;
always @(posedge clk)
m0122<=h012201;
always @(posedge clk)
m0123<=h012301;
always @(posedge clk)
m0124<=h012401;
always @(posedge clk)
m0125<=h012501;
always @(posedge clk)
m0126<=h012601;
always @(posedge clk)
m0127<=h012701;
always @(posedge clk)
m0128<=h012801;
always @(posedge clk)
m0129<=h012901;
always @(posedge clk)
m0130<=h013001;
always @(posedge clk)
m0131<=h013101;
always @(posedge clk)
m0132<=h013201;
always @(posedge clk)
m0133<=h013301;
always @(posedge clk)
m0134<=h013401;
always @(posedge clk)
m0135<=h013501;
always @(posedge clk)
m0136<=h013601;
always @(posedge clk)
m0137<=h013701;
always @(posedge clk)
m0138<=h013801;
always @(posedge clk)
m0139<=h013901;
always @(posedge clk)
m0140<=h014001;
always @(posedge clk)
m0141<=h014101;
always @(posedge clk)
m0142<=h014201;
always @(posedge clk)
m0143<=h014301;
always @(posedge clk)
m0144<=h014401;
always @(posedge clk)
m0145<=h014501;
always @(posedge clk)
m0146<=h014601;
always @(posedge clk)
m0147<=h014701;
always @(posedge clk)
m0148<=h014801;
always @(posedge clk)
m0149<=h014901;
always @(posedge clk)
m0150<=h015001;

always @(negedge clk)
q0121<=m0121;
always @(negedge clk)
q0122<=m0122;
always @(negedge clk)
q0123<=m0123;
always @(negedge clk)
q0124<=m0124;
always @(negedge clk)
q0125<=m0125;
always @(negedge clk)
q0126<=m0126;
always @(negedge clk)
q0127<=m0127;
always @(negedge clk)
q0128<=m0128;
always @(negedge clk)
q0129<=m0129;
always @(negedge clk)
q0130<=m0130;
always @(negedge clk)
q0131<=m0131;
always @(negedge clk)
q0132<=m0132;
always @(negedge clk)
q0133<=m0133;
always @(negedge clk)
q0134<=m0134;
always @(negedge clk)
q0135<=m0135;
always @(negedge clk)
q0136<=m0136;
always @(negedge clk)
q0137<=m0137;
always @(negedge clk)
q0138<=m0138;
always @(negedge clk)
q0139<=m0139;
always @(negedge clk)
q0140<=m0140;
always @(negedge clk)
q0141<=m0141;
always @(negedge clk)
q0142<=m0142;
always @(negedge clk)
q0143<=m0143;
always @(negedge clk)
q0144<=m0144;
always @(negedge clk)
q0145<=m0145;
always @(negedge clk)
q0146<=m0146;
always @(negedge clk)
q0147<=m0147;
always @(negedge clk)
q0148<=m0148;
always @(negedge clk)
q0149<=m0149;
always @(negedge clk)
q0150<=m0150;
//1
always @(posedge clk)
m0151<=a0181;
always @(posedge clk)
m0152<=a0182;
always @(posedge clk)
m0153<=a0183;
always @(posedge clk)
m0154<=a0184;
always @(posedge clk)
m0155<=a0185;
always @(posedge clk)
m0156<=a0186;
always @(posedge clk)
m0157<=a0187;
always @(posedge clk)
m0158<=a0188;
always @(posedge clk)
m0159<=a0189;
always @(posedge clk)
m0160<=a0190;
always @(posedge clk)
m0161<=a0191;
always @(posedge clk)
m0162<=a0192;
always @(posedge clk)
m0163<=a0193;
always @(posedge clk)
m0164<=a0194;
always @(posedge clk)
m0165<=a0195;
always @(posedge clk)
m0166<=a0196;
always @(posedge clk)
m0167<=a0197;
always @(posedge clk)
m0168<=a0198;
always @(posedge clk)
m0169<=a0199;
always @(posedge clk)
m0170<=a0200;
always @(posedge clk)
m0171<=a0201;
always @(posedge clk)
m0172<=a0202;
always @(posedge clk)
m0173<=a0203;
always @(posedge clk)
m0174<=a0204;
always @(posedge clk)
m0175<=a0205;
always @(posedge clk)
m0176<=a0206;
always @(posedge clk)
m0177<=a0207;
always @(posedge clk)
m0178<=a0208;
always @(posedge clk)
m0179<=a0209;
always @(posedge clk)
m0180<=a0210;

always @(negedge clk)
q0151<=m0151;
always @(negedge clk)
q0152<=m0152;
always @(negedge clk)
q0153<=m0153;
always @(negedge clk)
q0154<=m0154;
always @(negedge clk)
q0155<=m0155;
always @(negedge clk)
q0156<=m0156;
always @(negedge clk)
q0157<=m0157;
always @(negedge clk)
q0158<=m0158;
always @(negedge clk)
q0159<=m0159;
always @(negedge clk)
q0160<=m0160;
always @(negedge clk)
q0161<=m0161;
always @(negedge clk)
q0162<=m0162;
always @(negedge clk)
q0163<=m0163;
always @(negedge clk)
q0164<=m0164;
always @(negedge clk)
q0165<=m0165;
always @(negedge clk)
q0166<=m0166;
always @(negedge clk)
q0167<=m0167;
always @(negedge clk)
q0168<=m0168;
always @(negedge clk)
q0169<=m0169;
always @(negedge clk)
q0170<=m0170;
always @(negedge clk)
q0171<=m0171;
always @(negedge clk)
q0172<=m0172;
always @(negedge clk)
q0173<=m0173;
always @(negedge clk)
q0174<=m0174;
always @(negedge clk)
q0175<=m0175;
always @(negedge clk)
q0176<=m0176;
always @(negedge clk)
q0177<=m0177;
always @(negedge clk)
q0178<=m0178;
always @(negedge clk)
q0179<=m0179;
always @(negedge clk)
q0180<=m0180;

always @(posedge clk)
m0181<=h018101;
always @(posedge clk)
m0182<=h018201;
always @(posedge clk)
m0183<=h018301;
always @(posedge clk)
m0184<=h018401;
always @(posedge clk)
m0185<=h018501;
always @(posedge clk)
m0186<=h018601;
always @(posedge clk)
m0187<=h018701;
always @(posedge clk)
m0188<=h018801;
always @(posedge clk)
m0189<=h018901;
always @(posedge clk)
m0190<=h019001;
always @(posedge clk)
m0191<=h019101;
always @(posedge clk)
m0192<=h019201;
always @(posedge clk)
m0193<=h019301;
always @(posedge clk)
m0194<=h019401;
always @(posedge clk)
m0195<=h019501;
always @(posedge clk)
m0196<=h019601;
always @(posedge clk)
m0197<=h019701;
always @(posedge clk)
m0198<=h019801;
always @(posedge clk)
m0199<=h019901;
always @(posedge clk)
m0200<=h020001;
always @(posedge clk)
m0201<=h020101;
always @(posedge clk)
m0202<=h020201;
always @(posedge clk)
m0203<=h020301;
always @(posedge clk)
m0204<=h020401;
always @(posedge clk)
m0205<=h020501;
always @(posedge clk)
m0206<=h020601;
always @(posedge clk)
m0207<=h020701;
always @(posedge clk)
m0208<=h020801;
always @(posedge clk)
m0209<=h020901;
always @(posedge clk)
m0210<=h021001;

always @(negedge clk)
q0181<=m0181;
always @(negedge clk)
q0182<=m0182;
always @(negedge clk)
q0183<=m0183;
always @(negedge clk)
q0184<=m0184;
always @(negedge clk)
q0185<=m0185;
always @(negedge clk)
q0186<=m0186;
always @(negedge clk)
q0187<=m0187;
always @(negedge clk)
q0188<=m0188;
always @(negedge clk)
q0189<=m0189;
always @(negedge clk)
q0190<=m0190;
always @(negedge clk)
q0191<=m0191;
always @(negedge clk)
q0192<=m0192;
always @(negedge clk)
q0193<=m0193;
always @(negedge clk)
q0194<=m0194;
always @(negedge clk)
q0195<=m0195;
always @(negedge clk)
q0196<=m0196;
always @(negedge clk)
q0197<=m0197;
always @(negedge clk)
q0198<=m0198;
always @(negedge clk)
q0199<=m0199;
always @(negedge clk)
q0200<=m0200;
always @(negedge clk)
q0201<=m0201;
always @(negedge clk)
q0202<=m0202;
always @(negedge clk)
q0203<=m0203;
always @(negedge clk)
q0204<=m0204;
always @(negedge clk)
q0205<=m0205;
always @(negedge clk)
q0206<=m0206;
always @(negedge clk)
q0207<=m0207;
always @(negedge clk)
q0208<=m0208;
always @(negedge clk)
q0209<=m0209;
always @(negedge clk)
q0210<=m0210;
//2
always @(posedge clk)
m0211<=a0241;
always @(posedge clk)
m0212<=a0242;
always @(posedge clk)
m0213<=a0243;
always @(posedge clk)
m0214<=a0244;
always @(posedge clk)
m0215<=a0245;
always @(posedge clk)
m0216<=a0246;
always @(posedge clk)
m0217<=a0247;
always @(posedge clk)
m0218<=a0248;
always @(posedge clk)
m0219<=a0249;
always @(posedge clk)
m0220<=a0250;
always @(posedge clk)
m0221<=a0251;
always @(posedge clk)
m0222<=a0252;
always @(posedge clk)
m0223<=a0253;
always @(posedge clk)
m0224<=a0254;
always @(posedge clk)
m0225<=a0255;
always @(posedge clk)
m0226<=a0256;
always @(posedge clk)
m0227<=a0257;
always @(posedge clk)
m0228<=a0258;
always @(posedge clk)
m0229<=a0259;
always @(posedge clk)
m0230<=a0260;
always @(posedge clk)
m0231<=a0261;
always @(posedge clk)
m0232<=a0262;
always @(posedge clk)
m0233<=a0263;
always @(posedge clk)
m0234<=a0264;
always @(posedge clk)
m0235<=a0265;
always @(posedge clk)
m0236<=a0266;
always @(posedge clk)
m0237<=a0267;
always @(posedge clk)
m0238<=a0268;
always @(posedge clk)
m0239<=a0269;
always @(posedge clk)
m0240<=a0270;

always @(negedge clk)
q0211<=m0211;
always @(negedge clk)
q0212<=m0212;
always @(negedge clk)
q0213<=m0213;
always @(negedge clk)
q0214<=m0214;
always @(negedge clk)
q0215<=m0215;
always @(negedge clk)
q0216<=m0216;
always @(negedge clk)
q0217<=m0217;
always @(negedge clk)
q0218<=m0218;
always @(negedge clk)
q0219<=m0219;
always @(negedge clk)
q0220<=m0220;
always @(negedge clk)
q0221<=m0221;
always @(negedge clk)
q0222<=m0222;
always @(negedge clk)
q0223<=m0223;
always @(negedge clk)
q0224<=m0224;
always @(negedge clk)
q0225<=m0225;
always @(negedge clk)
q0226<=m0226;
always @(negedge clk)
q0227<=m0227;
always @(negedge clk)
q0228<=m0228;
always @(negedge clk)
q0229<=m0229;
always @(negedge clk)
q0230<=m0230;
always @(negedge clk)
q0231<=m0231;
always @(negedge clk)
q0232<=m0232;
always @(negedge clk)
q0233<=m0233;
always @(negedge clk)
q0234<=m0234;
always @(negedge clk)
q0235<=m0235;
always @(negedge clk)
q0236<=m0236;
always @(negedge clk)
q0237<=m0237;
always @(negedge clk)
q0238<=m0238;
always @(negedge clk)
q0239<=m0239;
always @(negedge clk)
q0240<=m0240;

always @(posedge clk)
m0241<=h024101;
always @(posedge clk)
m0242<=h024201;
always @(posedge clk)
m0243<=h024301;
always @(posedge clk)
m0244<=h024401;
always @(posedge clk)
m0245<=h024501;
always @(posedge clk)
m0246<=h024601;
always @(posedge clk)
m0247<=h024701;
always @(posedge clk)
m0248<=h024801;
always @(posedge clk)
m0249<=h024901;
always @(posedge clk)
m0250<=h025001;
always @(posedge clk)
m0251<=h025101;
always @(posedge clk)
m0252<=h025201;
always @(posedge clk)
m0253<=h025301;
always @(posedge clk)
m0254<=h025401;
always @(posedge clk)
m0255<=h025501;
always @(posedge clk)
m0256<=h025601;
always @(posedge clk)
m0257<=h025701;
always @(posedge clk)
m0258<=h025801;
always @(posedge clk)
m0259<=h025901;
always @(posedge clk)
m0260<=h026001;
always @(posedge clk)
m0261<=h026101;
always @(posedge clk)
m0262<=h026201;
always @(posedge clk)
m0263<=h026301;
always @(posedge clk)
m0264<=h026401;
always @(posedge clk)
m0265<=h026501;
always @(posedge clk)
m0266<=h026601;
always @(posedge clk)
m0267<=h026701;
always @(posedge clk)
m0268<=h026801;
always @(posedge clk)
m0269<=h026901;
always @(posedge clk)
m0270<=h027001;

always @(negedge clk)
q0241<=m0241;
always @(negedge clk)
q0242<=m0242;
always @(negedge clk)
q0243<=m0243;
always @(negedge clk)
q0244<=m0244;
always @(negedge clk)
q0245<=m0245;
always @(negedge clk)
q0246<=m0246;
always @(negedge clk)
q0247<=m0247;
always @(negedge clk)
q0248<=m0248;
always @(negedge clk)
q0249<=m0249;
always @(negedge clk)
q0250<=m0250;
always @(negedge clk)
q0251<=m0251;
always @(negedge clk)
q0252<=m0252;
always @(negedge clk)
q0253<=m0253;
always @(negedge clk)
q0254<=m0254;
always @(negedge clk)
q0255<=m0255;
always @(negedge clk)
q0256<=m0256;
always @(negedge clk)
q0257<=m0257;
always @(negedge clk)
q0258<=m0258;
always @(negedge clk)
q0259<=m0259;
always @(negedge clk)
q0260<=m0260;
always @(negedge clk)
q0261<=m0261;
always @(negedge clk)
q0262<=m0262;
always @(negedge clk)
q0263<=m0263;
always @(negedge clk)
q0264<=m0264;
always @(negedge clk)
q0265<=m0265;
always @(negedge clk)
q0266<=m0266;
always @(negedge clk)
q0267<=m0267;
always @(negedge clk)
q0268<=m0268;
always @(negedge clk)
q0269<=m0269;
always @(negedge clk)
q0270<=m0270;
//s
always @(posedge clk)
m0271<=a0301;
always @(posedge clk)
m0272<=a0302;
always @(posedge clk)
m0273<=a0303;
always @(posedge clk)
m0274<=a0304;
always @(posedge clk)
m0275<=a0305;
always @(posedge clk)
m0276<=a0306;
always @(posedge clk)
m0277<=a0307;
always @(posedge clk)
m0278<=a0308;
always @(posedge clk)
m0279<=a0309;
always @(posedge clk)
m0280<=a0310;
always @(posedge clk)
m0281<=a0311;
always @(posedge clk)
m0282<=a0312;
always @(posedge clk)
m0283<=a0313;
always @(posedge clk)
m0284<=a0314;
always @(posedge clk)
m0285<=a0315;
always @(posedge clk)
m0286<=a0316;
always @(posedge clk)
m0287<=a0317;
always @(posedge clk)
m0288<=a0318;
always @(posedge clk)
m0289<=a0319;
always @(posedge clk)
m0290<=a0320;
always @(posedge clk)
m0291<=a0321;
always @(posedge clk)
m0292<=a0322;
always @(posedge clk)
m0293<=a0323;
always @(posedge clk)
m0294<=a0324;
always @(posedge clk)
m0295<=a0325;
always @(posedge clk)
m0296<=a0326;
always @(posedge clk)
m0297<=a0327;
always @(posedge clk)
m0298<=a0328;
always @(posedge clk)
m0299<=a0329;
always @(posedge clk)
m0300<=a0330;

always @(negedge clk)
q0271<=m0271;
always @(negedge clk)
q0272<=m0272;
always @(negedge clk)
q0273<=m0273;
always @(negedge clk)
q0274<=m0274;
always @(negedge clk)
q0275<=m0275;
always @(negedge clk)
q0276<=m0276;
always @(negedge clk)
q0277<=m0277;
always @(negedge clk)
q0278<=m0278;
always @(negedge clk)
q0279<=m0279;
always @(negedge clk)
q0280<=m0280;
always @(negedge clk)
q0281<=m0281;
always @(negedge clk)
q0282<=m0282;
always @(negedge clk)
q0283<=m0283;
always @(negedge clk)
q0284<=m0284;
always @(negedge clk)
q0285<=m0285;
always @(negedge clk)
q0286<=m0286;
always @(negedge clk)
q0287<=m0287;
always @(negedge clk)
q0288<=m0288;
always @(negedge clk)
q0289<=m0289;
always @(negedge clk)
q0290<=m0290;
always @(negedge clk)
q0291<=m0291;
always @(negedge clk)
q0292<=m0292;
always @(negedge clk)
q0293<=m0293;
always @(negedge clk)
q0294<=m0294;
always @(negedge clk)
q0295<=m0295;
always @(negedge clk)
q0296<=m0296;
always @(negedge clk)
q0297<=m0297;
always @(negedge clk)
q0298<=m0298;
always @(negedge clk)
q0299<=m0299;
always @(negedge clk)
q0300<=m0300;

always @(posedge clk)
m0301<=h030101;
always @(posedge clk)
m0302<=h030201;
always @(posedge clk)
m0303<=h030301;
always @(posedge clk)
m0304<=h030401;
always @(posedge clk)
m0305<=h030501;
always @(posedge clk)
m0306<=h030601;
always @(posedge clk)
m0307<=h030701;
always @(posedge clk)
m0308<=h030801;
always @(posedge clk)
m0309<=h030901;
always @(posedge clk)
m0310<=h031001;
always @(posedge clk)
m0311<=h031101;
always @(posedge clk)
m0312<=h031201;
always @(posedge clk)
m0313<=h031301;
always @(posedge clk)
m0314<=h031401;
always @(posedge clk)
m0315<=h031501;
always @(posedge clk)
m0316<=h031601;
always @(posedge clk)
m0317<=h031701;
always @(posedge clk)
m0318<=h031801;
always @(posedge clk)
m0319<=h031901;
always @(posedge clk)
m0320<=h032001;
always @(posedge clk)
m0321<=h032101;
always @(posedge clk)
m0322<=h032201;
always @(posedge clk)
m0323<=h032301;
always @(posedge clk)
m0324<=h032401;
always @(posedge clk)
m0325<=h032501;
always @(posedge clk)
m0326<=h032601;
always @(posedge clk)
m0327<=h032701;
always @(posedge clk)
m0328<=h032801;
always @(posedge clk)
m0329<=h032901;
always @(posedge clk)
m0330<=h033001;

always @(negedge clk)
q0301<=m0301;
always @(negedge clk)
q0302<=m0302;
always @(negedge clk)
q0303<=m0303;
always @(negedge clk)
q0304<=m0304;
always @(negedge clk)
q0305<=m0305;
always @(negedge clk)
q0306<=m0306;
always @(negedge clk)
q0307<=m0307;
always @(negedge clk)
q0308<=m0308;
always @(negedge clk)
q0309<=m0309;
always @(negedge clk)
q0310<=m0310;
always @(negedge clk)
q0311<=m0311;
always @(negedge clk)
q0312<=m0312;
always @(negedge clk)
q0313<=m0313;
always @(negedge clk)
q0314<=m0314;
always @(negedge clk)
q0315<=m0315;
always @(negedge clk)
q0316<=m0316;
always @(negedge clk)
q0317<=m0317;
always @(negedge clk)
q0318<=m0318;
always @(negedge clk)
q0319<=m0319;
always @(negedge clk)
q0320<=m0320;
always @(negedge clk)
q0321<=m0321;
always @(negedge clk)
q0322<=m0322;
always @(negedge clk)
q0323<=m0323;
always @(negedge clk)
q0324<=m0324;
always @(negedge clk)
q0325<=m0325;
always @(negedge clk)
q0326<=m0326;
always @(negedge clk)
q0327<=m0327;
always @(negedge clk)
q0328<=m0328;
always @(negedge clk)
q0329<=m0329;
always @(negedge clk)
q0330<=m0330;
//so
always @(posedge clk)
m0331<=a0361;
always @(posedge clk)
m0332<=a0362;
always @(posedge clk)
m0333<=a0363;
always @(posedge clk)
m0334<=a0364;
always @(posedge clk)
m0335<=a0365;
always @(posedge clk)
m0336<=a0366;
always @(posedge clk)
m0337<=a0367;
always @(posedge clk)
m0338<=a0368;
always @(posedge clk)
m0339<=a0369;
always @(posedge clk)
m0340<=a0370;
always @(posedge clk)
m0341<=a0371;
always @(posedge clk)
m0342<=a0372;
always @(posedge clk)
m0343<=a0373;
always @(posedge clk)
m0344<=a0374;
always @(posedge clk)
m0345<=a0375;
always @(posedge clk)
m0346<=a0376;
always @(posedge clk)
m0347<=a0377;
always @(posedge clk)
m0348<=a0378;
always @(posedge clk)
m0349<=a0379;
always @(posedge clk)
m0350<=a0380;
always @(posedge clk)
m0351<=a0381;
always @(posedge clk)
m0352<=a0382;
always @(posedge clk)
m0353<=a0383;
always @(posedge clk)
m0354<=a0384;
always @(posedge clk)
m0355<=a0385;
always @(posedge clk)
m0356<=a0386;
always @(posedge clk)
m0357<=a0387;
always @(posedge clk)
m0358<=a0388;
always @(posedge clk)
m0359<=a0389;
always @(posedge clk)
m0360<=a0390;

always @(negedge clk)
q0331<=m0331;
always @(negedge clk)
q0332<=m0332;
always @(negedge clk)
q0333<=m0333;
always @(negedge clk)
q0334<=m0334;
always @(negedge clk)
q0335<=m0335;
always @(negedge clk)
q0336<=m0336;
always @(negedge clk)
q0337<=m0337;
always @(negedge clk)
q0338<=m0338;
always @(negedge clk)
q0339<=m0339;
always @(negedge clk)
q0340<=m0340;
always @(negedge clk)
q0341<=m0341;
always @(negedge clk)
q0342<=m0342;
always @(negedge clk)
q0343<=m0343;
always @(negedge clk)
q0344<=m0344;
always @(negedge clk)
q0345<=m0345;
always @(negedge clk)
q0346<=m0346;
always @(negedge clk)
q0347<=m0347;
always @(negedge clk)
q0348<=m0348;
always @(negedge clk)
q0349<=m0349;
always @(negedge clk)
q0350<=m0350;
always @(negedge clk)
q0351<=m0351;
always @(negedge clk)
q0352<=m0352;
always @(negedge clk)
q0353<=m0353;
always @(negedge clk)
q0354<=m0354;
always @(negedge clk)
q0355<=m0355;
always @(negedge clk)
q0356<=m0356;
always @(negedge clk)
q0357<=m0357;
always @(negedge clk)
q0358<=m0358;
always @(negedge clk)
q0359<=m0359;
always @(negedge clk)
q0360<=m0360;

always @(posedge clk)
m0361<=h036101;
always @(posedge clk)
m0362<=h036201;
always @(posedge clk)
m0363<=h036301;
always @(posedge clk)
m0364<=h036401;
always @(posedge clk)
m0365<=h036501;
always @(posedge clk)
m0366<=h036601;
always @(posedge clk)
m0367<=h036701;
always @(posedge clk)
m0368<=h036801;
always @(posedge clk)
m0369<=h036901;
always @(posedge clk)
m0370<=h037001;
always @(posedge clk)
m0371<=h037101;
always @(posedge clk)
m0372<=h037201;
always @(posedge clk)
m0373<=h037301;
always @(posedge clk)
m0374<=h037401;
always @(posedge clk)
m0375<=h037501;
always @(posedge clk)
m0376<=h037601;
always @(posedge clk)
m0377<=h037701;
always @(posedge clk)
m0378<=h037801;
always @(posedge clk)
m0379<=h037901;
always @(posedge clk)
m0380<=h038001;
always @(posedge clk)
m0381<=h038101;
always @(posedge clk)
m0382<=h038201;
always @(posedge clk)
m0383<=h038301;
always @(posedge clk)
m0384<=h038401;
always @(posedge clk)
m0385<=h038501;
always @(posedge clk)
m0386<=h038601;
always @(posedge clk)
m0387<=h038701;
always @(posedge clk)
m0388<=h038801;
always @(posedge clk)
m0389<=h038901;
always @(posedge clk)
m0390<=h039001;

always @(negedge clk)
q0361<=m0361;
always @(negedge clk)
q0362<=m0362;
always @(negedge clk)
q0363<=m0363;
always @(negedge clk)
q0364<=m0364;
always @(negedge clk)
q0365<=m0365;
always @(negedge clk)
q0366<=m0366;
always @(negedge clk)
q0367<=m0367;
always @(negedge clk)
q0368<=m0368;
always @(negedge clk)
q0369<=m0369;
always @(negedge clk)
q0370<=m0370;
always @(negedge clk)
q0371<=m0371;
always @(negedge clk)
q0372<=m0372;
always @(negedge clk)
q0373<=m0373;
always @(negedge clk)
q0374<=m0374;
always @(negedge clk)
q0375<=m0375;
always @(negedge clk)
q0376<=m0376;
always @(negedge clk)
q0377<=m0377;
always @(negedge clk)
q0378<=m0378;
always @(negedge clk)
q0379<=m0379;
always @(negedge clk)
q0380<=m0380;
always @(negedge clk)
q0381<=m0381;
always @(negedge clk)
q0382<=m0382;
always @(negedge clk)
q0383<=m0383;
always @(negedge clk)
q0384<=m0384;
always @(negedge clk)
q0385<=m0385;
always @(negedge clk)
q0386<=m0386;
always @(negedge clk)
q0387<=m0387;
always @(negedge clk)
q0388<=m0388;
always @(negedge clk)
q0389<=m0389;
always @(negedge clk)
q0390<=m0390;

always @(posedge clk)
m100_0<=h100_0;
always @(posedge clk)
m100_1<=h100_1;
always @(posedge clk)
m101_0<=h101_0;
always @(posedge clk)
m101_1<=h101_1;
always @(posedge clk)
m162_0<=h162_0;
always @(posedge clk)
m162_1<=h162_1;
always @(posedge clk)
m163_0<=h163_0;
always @(posedge clk)
m163_1<=h163_1;

always @(negedge clk)
q100_0<=m100_0;
always @(negedge clk)
q100_1<=m100_1;
always @(negedge clk)
q101_0<=m101_0;
always @(negedge clk)
q101_1<=m101_1;
always @(negedge clk)
q162_0<=m162_0;
always @(negedge clk)
q162_1<=m162_1;
always @(negedge clk)
q163_0<=m163_0;
always @(negedge clk)
q163_1<=m163_1;

always @(posedge clk)
m200_0<=h200_0;
always @(posedge clk)
m200_1<=h200_1;
always @(posedge clk)
m201_0<=h201_0;
always @(posedge clk)
m201_1<=h201_1;
always @(posedge clk)
m262_0<=h262_0;
always @(posedge clk)
m262_1<=h262_1;
always @(posedge clk)
m263_0<=h263_0;
always @(posedge clk)
m263_1<=h263_1;

always @(negedge clk)
q200_0<=m200_0;
always @(negedge clk)
q200_1<=m200_1;
always @(negedge clk)
q201_0<=m201_0;
always @(negedge clk)
q201_1<=m201_1;
always @(negedge clk)
q262_0<=m262_0;
always @(negedge clk)
q262_1<=m262_1;
always @(negedge clk)
q263_0<=m263_0;
always @(negedge clk)
q263_1<=m263_1;

always @(posedge clk)
m102_0<=h102_0;
always @(posedge clk)
m102_1<=h102_1;
always @(posedge clk)
m103_0<=h103_0;
always @(posedge clk)
m103_1<=h103_1;
always @(posedge clk)
m104_0<=h104_0;
always @(posedge clk)
m104_1<=h104_1;
always @(posedge clk)
m105_0<=h105_0;
always @(posedge clk)
m105_1<=h105_1;
always @(posedge clk)
m106_0<=h106_0;
always @(posedge clk)
m106_1<=h106_1;
always @(posedge clk)
m107_0<=h107_0;
always @(posedge clk)
m107_1<=h107_1;
always @(posedge clk)
m108_0<=h108_0;
always @(posedge clk)
m108_1<=h108_1;
always @(posedge clk)
m109_0<=h109_0;
always @(posedge clk)
m109_1<=h109_1;
always @(posedge clk)
m110_0<=h110_0;
always @(posedge clk)
m110_1<=h110_1;
always @(posedge clk)
m111_0<=h111_0;
always @(posedge clk)
m111_1<=h111_1;
always @(posedge clk)
m112_0<=h112_0;
always @(posedge clk)
m112_1<=h112_1;
always @(posedge clk)
m113_0<=h113_0;
always @(posedge clk)
m113_1<=h113_1;
always @(posedge clk)
m114_0<=h114_0;
always @(posedge clk)
m114_1<=h114_1;
always @(posedge clk)
m115_0<=h115_0;
always @(posedge clk)
m115_1<=h115_1;
always @(posedge clk)
m116_0<=h116_0;
always @(posedge clk)
m116_1<=h116_1;
always @(posedge clk)
m117_0<=h117_0;
always @(posedge clk)
m117_1<=h117_1;
always @(posedge clk)
m118_0<=h118_0;
always @(posedge clk)
m118_1<=h118_1;
always @(posedge clk)
m119_0<=h119_0;
always @(posedge clk)
m119_1<=h119_1;
always @(posedge clk)
m120_0<=h120_0;
always @(posedge clk)
m120_1<=h120_1;
always @(posedge clk)
m121_0<=h121_0;
always @(posedge clk)
m121_1<=h121_1;
always @(posedge clk)
m122_0<=h122_0;
always @(posedge clk)
m122_1<=h122_1;
always @(posedge clk)
m123_0<=h123_0;
always @(posedge clk)
m123_1<=h123_1;
always @(posedge clk)
m124_0<=h124_0;
always @(posedge clk)
m124_1<=h124_1;
always @(posedge clk)
m125_0<=h125_0;
always @(posedge clk)
m125_1<=h125_1;
always @(posedge clk)
m126_0<=h126_0;
always @(posedge clk)
m126_1<=h126_1;
always @(posedge clk)
m127_0<=h127_0;
always @(posedge clk)
m127_1<=h127_1;
always @(posedge clk)
m128_0<=h128_0;
always @(posedge clk)
m128_1<=h128_1;
always @(posedge clk)
m129_0<=h129_0;
always @(posedge clk)
m129_1<=h129_1;
always @(posedge clk)
m130_0<=h130_0;
always @(posedge clk)
m130_1<=h130_1;
always @(posedge clk)
m131_0<=h131_0;
always @(posedge clk)
m131_1<=h131_1;
always @(posedge clk)
m132_0<=h132_0;
always @(posedge clk)
m132_1<=h132_1;
always @(posedge clk)
m133_0<=h133_0;
always @(posedge clk)
m133_1<=h133_1;
always @(posedge clk)
m134_0<=h134_0;
always @(posedge clk)
m134_1<=h134_1;
always @(posedge clk)
m135_0<=h135_0;
always @(posedge clk)
m135_1<=h135_1;
always @(posedge clk)
m136_0<=h136_0;
always @(posedge clk)
m136_1<=h136_1;
always @(posedge clk)
m137_0<=h137_0;
always @(posedge clk)
m137_1<=h137_1;
always @(posedge clk)
m138_0<=h138_0;
always @(posedge clk)
m138_1<=h138_1;
always @(posedge clk)
m139_0<=h139_0;
always @(posedge clk)
m139_1<=h139_1;
always @(posedge clk)
m140_0<=h140_0;
always @(posedge clk)
m140_1<=h140_1;
always @(posedge clk)
m141_0<=h141_0;
always @(posedge clk)
m141_1<=h141_1;
always @(posedge clk)
m142_0<=h142_0;
always @(posedge clk)
m142_1<=h142_1;
always @(posedge clk)
m143_0<=h143_0;
always @(posedge clk)
m143_1<=h143_1;
always @(posedge clk)
m144_0<=h144_0;
always @(posedge clk)
m144_1<=h144_1;
always @(posedge clk)
m145_0<=h145_0;
always @(posedge clk)
m145_1<=h145_1;
always @(posedge clk)
m146_0<=h146_0;
always @(posedge clk)
m146_1<=h146_1;
always @(posedge clk)
m147_0<=h147_0;
always @(posedge clk)
m147_1<=h147_1;
always @(posedge clk)
m148_0<=h148_0;
always @(posedge clk)
m148_1<=h148_1;
always @(posedge clk)
m149_0<=h149_0;
always @(posedge clk)
m149_1<=h149_1;
always @(posedge clk)
m150_0<=h150_0;
always @(posedge clk)
m150_1<=h150_1;
always @(posedge clk)
m151_0<=h151_0;
always @(posedge clk)
m151_1<=h151_1;
always @(posedge clk)
m152_0<=h152_0;
always @(posedge clk)
m152_1<=h152_1;
always @(posedge clk)
m153_0<=h153_0;
always @(posedge clk)
m153_1<=h153_1;
always @(posedge clk)
m154_0<=h154_0;
always @(posedge clk)
m154_1<=h154_1;
always @(posedge clk)
m155_0<=h155_0;
always @(posedge clk)
m155_1<=h155_1;
always @(posedge clk)
m156_0<=h156_0;
always @(posedge clk)
m156_1<=h156_1;
always @(posedge clk)
m157_0<=h157_0;
always @(posedge clk)
m157_1<=h157_1;
always @(posedge clk)
m158_0<=h158_0;
always @(posedge clk)
m158_1<=h158_1;
always @(posedge clk)
m159_0<=h159_0;
always @(posedge clk)
m159_1<=h159_1;
always @(posedge clk)
m160_0<=h160_0;
always @(posedge clk)
m160_1<=h160_1;
always @(posedge clk)
m161_0<=h161_0;
always @(posedge clk)
m161_1<=h161_1;

always @(negedge clk)
q102_0<=m102_0;
always @(negedge clk)
q102_1<=m102_1;
always @(negedge clk)
q103_0<=m103_0;
always @(negedge clk)
q103_1<=m103_1;
always @(negedge clk)
q104_0<=m104_0;
always @(negedge clk)
q104_1<=m104_1;
always @(negedge clk)
q105_0<=m105_0;
always @(negedge clk)
q105_1<=m105_1;
always @(negedge clk)
q106_0<=m106_0;
always @(negedge clk)
q106_1<=m106_1;
always @(negedge clk)
q107_0<=m107_0;
always @(negedge clk)
q107_1<=m107_1;
always @(negedge clk)
q108_0<=m108_0;
always @(negedge clk)
q108_1<=m108_1;
always @(negedge clk)
q109_0<=m109_0;
always @(negedge clk)
q109_1<=m109_1;
always @(negedge clk)
q110_0<=m110_0;
always @(negedge clk)
q110_1<=m110_1;
always @(negedge clk)
q111_0<=m111_0;
always @(negedge clk)
q111_1<=m111_1;
always @(negedge clk)
q112_0<=m112_0;
always @(negedge clk)
q112_1<=m112_1;
always @(negedge clk)
q113_0<=m113_0;
always @(negedge clk)
q113_1<=m113_1;
always @(negedge clk)
q114_0<=m114_0;
always @(negedge clk)
q114_1<=m114_1;
always @(negedge clk)
q115_0<=m115_0;
always @(negedge clk)
q115_1<=m115_1;
always @(negedge clk)
q116_0<=m116_0;
always @(negedge clk)
q116_1<=m116_1;
always @(negedge clk)
q117_0<=m117_0;
always @(negedge clk)
q117_1<=m117_1;
always @(negedge clk)
q118_0<=m118_0;
always @(negedge clk)
q118_1<=m118_1;
always @(negedge clk)
q119_0<=m119_0;
always @(negedge clk)
q119_1<=m119_1;
always @(negedge clk)
q120_0<=m120_0;
always @(negedge clk)
q120_1<=m120_1;
always @(negedge clk)
q121_0<=m121_0;
always @(negedge clk)
q121_1<=m121_1;
always @(negedge clk)
q122_0<=m122_0;
always @(negedge clk)
q122_1<=m122_1;
always @(negedge clk)
q123_0<=m123_0;
always @(negedge clk)
q123_1<=m123_1;
always @(negedge clk)
q124_0<=m124_0;
always @(negedge clk)
q124_1<=m124_1;
always @(negedge clk)
q125_0<=m125_0;
always @(negedge clk)
q125_1<=m125_1;
always @(negedge clk)
q126_0<=m126_0;
always @(negedge clk)
q126_1<=m126_1;
always @(negedge clk)
q127_0<=m127_0;
always @(negedge clk)
q127_1<=m127_1;
always @(negedge clk)
q128_0<=m128_0;
always @(negedge clk)
q128_1<=m128_1;
always @(negedge clk)
q129_0<=m129_0;
always @(negedge clk)
q129_1<=m129_1;
always @(negedge clk)
q130_0<=m130_0;
always @(negedge clk)
q130_1<=m130_1;
always @(negedge clk)
q131_0<=m131_0;
always @(negedge clk)
q131_1<=m131_1;
always @(negedge clk)
q132_0<=m132_0;
always @(negedge clk)
q132_1<=m132_1;
always @(negedge clk)
q133_0<=m133_0;
always @(negedge clk)
q133_1<=m133_1;
always @(negedge clk)
q134_0<=m134_0;
always @(negedge clk)
q134_1<=m134_1;
always @(negedge clk)
q135_0<=m135_0;
always @(negedge clk)
q135_1<=m135_1;
always @(negedge clk)
q136_0<=m136_0;
always @(negedge clk)
q136_1<=m136_1;
always @(negedge clk)
q137_0<=m137_0;
always @(negedge clk)
q137_1<=m137_1;
always @(negedge clk)
q138_0<=m138_0;
always @(negedge clk)
q138_1<=m138_1;
always @(negedge clk)
q139_0<=m139_0;
always @(negedge clk)
q139_1<=m139_1;
always @(negedge clk)
q140_0<=m140_0;
always @(negedge clk)
q140_1<=m140_1;
always @(negedge clk)
q141_0<=m141_0;
always @(negedge clk)
q141_1<=m141_1;
always @(negedge clk)
q142_0<=m142_0;
always @(negedge clk)
q142_1<=m142_1;
always @(negedge clk)
q143_0<=m143_0;
always @(negedge clk)
q143_1<=m143_1;
always @(negedge clk)
q144_0<=m144_0;
always @(negedge clk)
q144_1<=m144_1;
always @(negedge clk)
q145_0<=m145_0;
always @(negedge clk)
q145_1<=m145_1;
always @(negedge clk)
q146_0<=m146_0;
always @(negedge clk)
q146_1<=m146_1;
always @(negedge clk)
q147_0<=m147_0;
always @(negedge clk)
q147_1<=m147_1;
always @(negedge clk)
q148_0<=m148_0;
always @(negedge clk)
q148_1<=m148_1;
always @(negedge clk)
q149_0<=m149_0;
always @(negedge clk)
q149_1<=m149_1;
always @(negedge clk)
q150_0<=m150_0;
always @(negedge clk)
q150_1<=m150_1;
always @(negedge clk)
q151_0<=m151_0;
always @(negedge clk)
q151_1<=m151_1;
always @(negedge clk)
q152_0<=m152_0;
always @(negedge clk)
q152_1<=m152_1;
always @(negedge clk)
q153_0<=m153_0;
always @(negedge clk)
q153_1<=m153_1;
always @(negedge clk)
q154_0<=m154_0;
always @(negedge clk)
q154_1<=m154_1;
always @(negedge clk)
q155_0<=m155_0;
always @(negedge clk)
q155_1<=m155_1;
always @(negedge clk)
q156_0<=m156_0;
always @(negedge clk)
q156_1<=m156_1;
always @(negedge clk)
q157_0<=m157_0;
always @(negedge clk)
q157_1<=m157_1;
always @(negedge clk)
q158_0<=m158_0;
always @(negedge clk)
q158_1<=m158_1;
always @(negedge clk)
q159_0<=m159_0;
always @(negedge clk)
q159_1<=m159_1;
always @(negedge clk)
q160_0<=m160_0;
always @(negedge clk)
q160_1<=m160_1;
always @(negedge clk)
q161_0<=m161_0;
always @(negedge clk)
q161_1<=m161_1;

always @(posedge clk)
m202_0<=h202_0;
always @(posedge clk)
m202_1<=h202_1;
always @(posedge clk)
m203_0<=h203_0;
always @(posedge clk)
m203_1<=h203_1;
always @(posedge clk)
m204_0<=h204_0;
always @(posedge clk)
m204_1<=h204_1;
always @(posedge clk)
m205_0<=h205_0;
always @(posedge clk)
m205_1<=h205_1;
always @(posedge clk)
m206_0<=h206_0;
always @(posedge clk)
m206_1<=h206_1;
always @(posedge clk)
m207_0<=h207_0;
always @(posedge clk)
m207_1<=h207_1;
always @(posedge clk)
m208_0<=h208_0;
always @(posedge clk)
m208_1<=h208_1;
always @(posedge clk)
m209_0<=h209_0;
always @(posedge clk)
m209_1<=h209_1;
always @(posedge clk)
m210_0<=h210_0;
always @(posedge clk)
m210_1<=h210_1;
always @(posedge clk)
m211_0<=h211_0;
always @(posedge clk)
m211_1<=h211_1;
always @(posedge clk)
m212_0<=h212_0;
always @(posedge clk)
m212_1<=h212_1;
always @(posedge clk)
m213_0<=h213_0;
always @(posedge clk)
m213_1<=h213_1;
always @(posedge clk)
m214_0<=h214_0;
always @(posedge clk)
m214_1<=h214_1;
always @(posedge clk)
m215_0<=h215_0;
always @(posedge clk)
m215_1<=h215_1;
always @(posedge clk)
m216_0<=h216_0;
always @(posedge clk)
m216_1<=h216_1;
always @(posedge clk)
m217_0<=h217_0;
always @(posedge clk)
m217_1<=h217_1;
always @(posedge clk)
m218_0<=h218_0;
always @(posedge clk)
m218_1<=h218_1;
always @(posedge clk)
m219_0<=h219_0;
always @(posedge clk)
m219_1<=h219_1;
always @(posedge clk)
m220_0<=h220_0;
always @(posedge clk)
m220_1<=h220_1;
always @(posedge clk)
m221_0<=h221_0;
always @(posedge clk)
m221_1<=h221_1;
always @(posedge clk)
m222_0<=h222_0;
always @(posedge clk)
m222_1<=h222_1;
always @(posedge clk)
m223_0<=h223_0;
always @(posedge clk)
m223_1<=h223_1;
always @(posedge clk)
m224_0<=h224_0;
always @(posedge clk)
m224_1<=h224_1;
always @(posedge clk)
m225_0<=h225_0;
always @(posedge clk)
m225_1<=h225_1;
always @(posedge clk)
m226_0<=h226_0;
always @(posedge clk)
m226_1<=h226_1;
always @(posedge clk)
m227_0<=h227_0;
always @(posedge clk)
m227_1<=h227_1;
always @(posedge clk)
m228_0<=h228_0;
always @(posedge clk)
m228_1<=h228_1;
always @(posedge clk)
m229_0<=h229_0;
always @(posedge clk)
m229_1<=h229_1;
always @(posedge clk)
m230_0<=h230_0;
always @(posedge clk)
m230_1<=h230_1;
always @(posedge clk)
m231_0<=h231_0;
always @(posedge clk)
m231_1<=h231_1;
always @(posedge clk)
m232_0<=h232_0;
always @(posedge clk)
m232_1<=h232_1;
always @(posedge clk)
m233_0<=h233_0;
always @(posedge clk)
m233_1<=h233_1;
always @(posedge clk)
m234_0<=h234_0;
always @(posedge clk)
m234_1<=h234_1;
always @(posedge clk)
m235_0<=h235_0;
always @(posedge clk)
m235_1<=h235_1;
always @(posedge clk)
m236_0<=h236_0;
always @(posedge clk)
m236_1<=h236_1;
always @(posedge clk)
m237_0<=h237_0;
always @(posedge clk)
m237_1<=h237_1;
always @(posedge clk)
m238_0<=h238_0;
always @(posedge clk)
m238_1<=h238_1;
always @(posedge clk)
m239_0<=h239_0;
always @(posedge clk)
m239_1<=h239_1;
always @(posedge clk)
m240_0<=h240_0;
always @(posedge clk)
m240_1<=h240_1;
always @(posedge clk)
m241_0<=h241_0;
always @(posedge clk)
m241_1<=h241_1;
always @(posedge clk)
m242_0<=h242_0;
always @(posedge clk)
m242_1<=h242_1;
always @(posedge clk)
m243_0<=h243_0;
always @(posedge clk)
m243_1<=h243_1;
always @(posedge clk)
m244_0<=h244_0;
always @(posedge clk)
m244_1<=h244_1;
always @(posedge clk)
m245_0<=h245_0;
always @(posedge clk)
m245_1<=h245_1;
always @(posedge clk)
m246_0<=h246_0;
always @(posedge clk)
m246_1<=h246_1;
always @(posedge clk)
m247_0<=h247_0;
always @(posedge clk)
m247_1<=h247_1;
always @(posedge clk)
m248_0<=h248_0;
always @(posedge clk)
m248_1<=h248_1;
always @(posedge clk)
m249_0<=h249_0;
always @(posedge clk)
m249_1<=h249_1;
always @(posedge clk)
m250_0<=h250_0;
always @(posedge clk)
m250_1<=h250_1;
always @(posedge clk)
m251_0<=h251_0;
always @(posedge clk)
m251_1<=h251_1;
always @(posedge clk)
m252_0<=h252_0;
always @(posedge clk)
m252_1<=h252_1;
always @(posedge clk)
m253_0<=h253_0;
always @(posedge clk)
m253_1<=h253_1;
always @(posedge clk)
m254_0<=h254_0;
always @(posedge clk)
m254_1<=h254_1;
always @(posedge clk)
m255_0<=h255_0;
always @(posedge clk)
m255_1<=h255_1;
always @(posedge clk)
m256_0<=h256_0;
always @(posedge clk)
m256_1<=h256_1;
always @(posedge clk)
m257_0<=h257_0;
always @(posedge clk)
m257_1<=h257_1;
always @(posedge clk)
m258_0<=h258_0;
always @(posedge clk)
m258_1<=h258_1;
always @(posedge clk)
m259_0<=h259_0;
always @(posedge clk)
m259_1<=h259_1;
always @(posedge clk)
m260_0<=h260_0;
always @(posedge clk)
m260_1<=h260_1;
always @(posedge clk)
m261_0<=h261_0;
always @(posedge clk)
m261_1<=h261_1;

always @(negedge clk)
q202_0<=m202_0;
always @(negedge clk)
q202_1<=m202_1;
always @(negedge clk)
q203_0<=m203_0;
always @(negedge clk)
q203_1<=m203_1;
always @(negedge clk)
q204_0<=m204_0;
always @(negedge clk)
q204_1<=m204_1;
always @(negedge clk)
q205_0<=m205_0;
always @(negedge clk)
q205_1<=m205_1;
always @(negedge clk)
q206_0<=m206_0;
always @(negedge clk)
q206_1<=m206_1;
always @(negedge clk)
q207_0<=m207_0;
always @(negedge clk)
q207_1<=m207_1;
always @(negedge clk)
q208_0<=m208_0;
always @(negedge clk)
q208_1<=m208_1;
always @(negedge clk)
q209_0<=m209_0;
always @(negedge clk)
q209_1<=m209_1;
always @(negedge clk)
q210_0<=m210_0;
always @(negedge clk)
q210_1<=m210_1;
always @(negedge clk)
q211_0<=m211_0;
always @(negedge clk)
q211_1<=m211_1;
always @(negedge clk)
q212_0<=m212_0;
always @(negedge clk)
q212_1<=m212_1;
always @(negedge clk)
q213_0<=m213_0;
always @(negedge clk)
q213_1<=m213_1;
always @(negedge clk)
q214_0<=m214_0;
always @(negedge clk)
q214_1<=m214_1;
always @(negedge clk)
q215_0<=m215_0;
always @(negedge clk)
q215_1<=m215_1;
always @(negedge clk)
q216_0<=m216_0;
always @(negedge clk)
q216_1<=m216_1;
always @(negedge clk)
q217_0<=m217_0;
always @(negedge clk)
q217_1<=m217_1;
always @(negedge clk)
q218_0<=m218_0;
always @(negedge clk)
q218_1<=m218_1;
always @(negedge clk)
q219_0<=m219_0;
always @(negedge clk)
q219_1<=m219_1;
always @(negedge clk)
q220_0<=m220_0;
always @(negedge clk)
q220_1<=m220_1;
always @(negedge clk)
q221_0<=m221_0;
always @(negedge clk)
q221_1<=m221_1;
always @(negedge clk)
q222_0<=m222_0;
always @(negedge clk)
q222_1<=m222_1;
always @(negedge clk)
q223_0<=m223_0;
always @(negedge clk)
q223_1<=m223_1;
always @(negedge clk)
q224_0<=m224_0;
always @(negedge clk)
q224_1<=m224_1;
always @(negedge clk)
q225_0<=m225_0;
always @(negedge clk)
q225_1<=m225_1;
always @(negedge clk)
q226_0<=m226_0;
always @(negedge clk)
q226_1<=m226_1;
always @(negedge clk)
q227_0<=m227_0;
always @(negedge clk)
q227_1<=m227_1;
always @(negedge clk)
q228_0<=m228_0;
always @(negedge clk)
q228_1<=m228_1;
always @(negedge clk)
q229_0<=m229_0;
always @(negedge clk)
q229_1<=m229_1;
always @(negedge clk)
q230_0<=m230_0;
always @(negedge clk)
q230_1<=m230_1;
always @(negedge clk)
q231_0<=m231_0;
always @(negedge clk)
q231_1<=m231_1;
always @(negedge clk)
q232_0<=m232_0;
always @(negedge clk)
q232_1<=m232_1;
always @(negedge clk)
q233_0<=m233_0;
always @(negedge clk)
q233_1<=m233_1;
always @(negedge clk)
q234_0<=m234_0;
always @(negedge clk)
q234_1<=m234_1;
always @(negedge clk)
q235_0<=m235_0;
always @(negedge clk)
q235_1<=m235_1;
always @(negedge clk)
q236_0<=m236_0;
always @(negedge clk)
q236_1<=m236_1;
always @(negedge clk)
q237_0<=m237_0;
always @(negedge clk)
q237_1<=m237_1;
always @(negedge clk)
q238_0<=m238_0;
always @(negedge clk)
q238_1<=m238_1;
always @(negedge clk)
q239_0<=m239_0;
always @(negedge clk)
q239_1<=m239_1;
always @(negedge clk)
q240_0<=m240_0;
always @(negedge clk)
q240_1<=m240_1;
always @(negedge clk)
q241_0<=m241_0;
always @(negedge clk)
q241_1<=m241_1;
always @(negedge clk)
q242_0<=m242_0;
always @(negedge clk)
q242_1<=m242_1;
always @(negedge clk)
q243_0<=m243_0;
always @(negedge clk)
q243_1<=m243_1;
always @(negedge clk)
q244_0<=m244_0;
always @(negedge clk)
q244_1<=m244_1;
always @(negedge clk)
q245_0<=m245_0;
always @(negedge clk)
q245_1<=m245_1;
always @(negedge clk)
q246_0<=m246_0;
always @(negedge clk)
q246_1<=m246_1;
always @(negedge clk)
q247_0<=m247_0;
always @(negedge clk)
q247_1<=m247_1;
always @(negedge clk)
q248_0<=m248_0;
always @(negedge clk)
q248_1<=m248_1;
always @(negedge clk)
q249_0<=m249_0;
always @(negedge clk)
q249_1<=m249_1;
always @(negedge clk)
q250_0<=m250_0;
always @(negedge clk)
q250_1<=m250_1;
always @(negedge clk)
q251_0<=m251_0;
always @(negedge clk)
q251_1<=m251_1;
always @(negedge clk)
q252_0<=m252_0;
always @(negedge clk)
q252_1<=m252_1;
always @(negedge clk)
q253_0<=m253_0;
always @(negedge clk)
q253_1<=m253_1;
always @(negedge clk)
q254_0<=m254_0;
always @(negedge clk)
q254_1<=m254_1;
always @(negedge clk)
q255_0<=m255_0;
always @(negedge clk)
q255_1<=m255_1;
always @(negedge clk)
q256_0<=m256_0;
always @(negedge clk)
q256_1<=m256_1;
always @(negedge clk)
q257_0<=m257_0;
always @(negedge clk)
q257_1<=m257_1;
always @(negedge clk)
q258_0<=m258_0;
always @(negedge clk)
q258_1<=m258_1;
always @(negedge clk)
q259_0<=m259_0;
always @(negedge clk)
q259_1<=m259_1;
always @(negedge clk)
q260_0<=m260_0;
always @(negedge clk)
q260_1<=m260_1;
always @(negedge clk)
q261_0<=m261_0;
always @(negedge clk)
q261_1<=m261_1;
/*
always @(posedge clk)
m1000_0<=h1000_0;
always @(posedge clk)
m1000_1<=h1000_1;
always @(posedge clk)
m1001_0<=h1001_0;
always @(posedge clk)
m1001_1<=h1001_1;
always @(posedge clk)
m1010_0<=h1010_0;
always @(posedge clk)
m1010_1<=h1010_1;
always @(posedge clk)
m1011_0<=h1011_0;
always @(posedge clk)
m1011_1<=h1011_1;
always @(posedge clk)
m1100_0<=h1100_0;
always @(posedge clk)
m1100_1<=h1100_1;
always @(posedge clk)
m1101_0<=h1101_0;
always @(posedge clk)
m1101_1<=h1101_1;
always @(posedge clk)
m1110_0<=h1110_0;
always @(posedge clk)
m1110_1<=h1110_1;
always @(posedge clk)
m1111_0<=h1111_0;
always @(posedge clk)
m1111_1<=h1111_1;

always @(negedge clk)
q1000_0<=m1000_0;
always @(negedge clk)
q1000_1<=m1000_1;
always @(negedge clk)
q1001_0<=m1001_0;
always @(negedge clk)
q1001_1<=m1001_1;
always @(negedge clk)
q1010_0<=m1010_0;
always @(negedge clk)
q1010_1<=m1010_1;
always @(negedge clk)
q1011_0<=m1011_0;
always @(negedge clk)
q1011_1<=m1011_1;
always @(negedge clk)
q1100_0<=m1100_0;
always @(negedge clk)
q1100_1<=m1100_1;
always @(negedge clk)
q1101_0<=m1101_0;
always @(negedge clk)
q1101_1<=m1101_1;
always @(negedge clk)
q1110_0<=m1110_0;
always @(negedge clk)
q1110_1<=m1110_1;
always @(negedge clk)
q1111_0<=m1111_0;
always @(negedge clk)
q1111_1<=m1111_1;

always @(posedge clk)
m2000_0<=h2000_0;
always @(posedge clk)
m2000_1<=h2000_1;
always @(posedge clk)
m2001_0<=h2001_0;
always @(posedge clk)
m2001_1<=h2001_1;
always @(posedge clk)
m2010_0<=h2010_0;
always @(posedge clk)
m2010_1<=h2010_1;
always @(posedge clk)
m2011_0<=h2011_0;
always @(posedge clk)
m2011_1<=h2011_1;
always @(posedge clk)
m2100_0<=h2100_0;
always @(posedge clk)
m2100_1<=h2100_1;
always @(posedge clk)
m2101_0<=h2101_0;
always @(posedge clk)
m2101_1<=h2101_1;
always @(posedge clk)
m2110_0<=h2110_0;
always @(posedge clk)
m2110_1<=h2110_1;
always @(posedge clk)
m2111_0<=h2111_0;
always @(posedge clk)
m2111_1<=h2111_1;

always @(negedge clk)
q2000_0<=m2000_0;
always @(negedge clk)
q2000_1<=m2000_1;
always @(negedge clk)
q2001_0<=m2001_0;
always @(negedge clk)
q2001_1<=m2001_1;
always @(negedge clk)
q2010_0<=m2010_0;
always @(negedge clk)
q2010_1<=m2010_1;
always @(negedge clk)
q2011_0<=m2011_0;
always @(negedge clk)
q2011_1<=m2011_1;
always @(negedge clk)
q2100_0<=m2100_0;
always @(negedge clk)
q2100_1<=m2100_1;
always @(negedge clk)
q2101_0<=m2101_0;
always @(negedge clk)
q2101_1<=m2101_1;
always @(negedge clk)
q2110_0<=m2110_0;
always @(negedge clk)
q2110_1<=m2110_1;
always @(negedge clk)
q2111_0<=m2111_0;
always @(negedge clk)
q2111_1<=m2111_1;
*/
always @(posedge clk)
m00_0<=h00_0;
always @(posedge clk)
m00_1<=h00_1;
always @(posedge clk)
m01_0<=h01_0;
always @(posedge clk)
m01_1<=h01_1;
always @(posedge clk)
m10_0<=h10_0;
always @(posedge clk)
m10_1<=h10_1;
always @(posedge clk)
m11_0<=h11_0;
always @(posedge clk)
m11_1<=h11_1;

always @(negedge clk)
q00_0<=m00_0;
always @(negedge clk)
q00_1<=m00_1;
always @(negedge clk)
q01_0<=m01_0;
always @(negedge clk)
q01_1<=m01_1;
always @(negedge clk)
q10_0<=m10_0;
always @(negedge clk)
q10_1<=m10_1;
always @(negedge clk)
q11_0<=m11_0;
always @(negedge clk)
q11_1<=m11_1;

always @(posedge clk)
ms_0<=hs_0;
always @(posedge clk)
ms_1<=hs_1;

always @(negedge clk)
qs_0<=ms_0;
always @(negedge clk)
qs_1<=ms_1;

always @(posedge clk)
mso_0<=hso_0;
always @(posedge clk)
mso_1<=hso_1;

always @(negedge clk)
qso_0<=mso_0;
always @(negedge clk)
qso_1<=mso_1;

always @(posedge clk)
m29_0<=h29_0;
always @(posedge clk)
m29_1<=h29_1;
always @(posedge clk)
m30_0<=h30_0;
always @(posedge clk)
m30_1<=h30_1;
always @(posedge clk)
m31_0<=h31_0;
always @(posedge clk)
m31_1<=h31_1;
always @(posedge clk)
m32_0<=h32_0;
always @(posedge clk)
m32_1<=h32_1;
always @(posedge clk)
m33_0<=h33_0;
always @(posedge clk)
m33_1<=h33_1;
always @(posedge clk)
m34_0<=h34_0;
always @(posedge clk)
m34_1<=h34_1;
always @(posedge clk)
m35_0<=h35_0;
always @(posedge clk)
m35_1<=h35_1;
always @(posedge clk)
m36_0<=h36_0;
always @(posedge clk)
m36_1<=h36_1;
always @(posedge clk)
m37_0<=h37_0;
always @(posedge clk)
m37_1<=h37_1;
always @(posedge clk)
m38_0<=h38_0;
always @(posedge clk)
m38_1<=h38_1;
always @(posedge clk)
m39_0<=h39_0;
always @(posedge clk)
m39_1<=h39_1;
always @(posedge clk)
m40_0<=h40_0;
always @(posedge clk)
m40_1<=h40_1;
always @(posedge clk)
m41_0<=h41_0;
always @(posedge clk)
m41_1<=h41_1;
always @(posedge clk)
m42_0<=h42_0;
always @(posedge clk)
m42_1<=h42_1;
always @(posedge clk)
m43_0<=h43_0;
always @(posedge clk)
m43_1<=h43_1;
always @(posedge clk)
m44_0<=h44_0;
always @(posedge clk)
m44_1<=h44_1;
always @(posedge clk)
m45_0<=h45_0;
always @(posedge clk)
m45_1<=h45_1;
always @(posedge clk)
m46_0<=h46_0;
always @(posedge clk)
m46_1<=h46_1;
always @(posedge clk)
m47_0<=h47_0;
always @(posedge clk)
m47_1<=h47_1;
always @(posedge clk)
m48_0<=h48_0;
always @(posedge clk)
m48_1<=h48_1;
always @(posedge clk)
m49_0<=h49_0;
always @(posedge clk)
m49_1<=h49_1;
always @(posedge clk)
m50_0<=h50_0;
always @(posedge clk)
m50_1<=h50_1;

always @(negedge clk)
q29_0<=m29_0;
always @(negedge clk)
q29_1<=m29_1;
always @(negedge clk)
q30_0<=m30_0;
always @(negedge clk)
q30_1<=m30_1;
always @(negedge clk)
q31_0<=m31_0;
always @(negedge clk)
q31_1<=m31_1;
always @(negedge clk)
q32_0<=m32_0;
always @(negedge clk)
q32_1<=m32_1;
always @(negedge clk)
q33_0<=m33_0;
always @(negedge clk)
q33_1<=m33_1;
always @(negedge clk)
q34_0<=m34_0;
always @(negedge clk)
q34_1<=m34_1;
always @(negedge clk)
q35_0<=m35_0;
always @(negedge clk)
q35_1<=m35_1;
always @(negedge clk)
q36_0<=m36_0;
always @(negedge clk)
q36_1<=m36_1;
always @(negedge clk)
q37_0<=m37_0;
always @(negedge clk)
q37_1<=m37_1;
always @(negedge clk)
q38_0<=m38_0;
always @(negedge clk)
q38_1<=m38_1;
always @(negedge clk)
q39_0<=m39_0;
always @(negedge clk)
q39_1<=m39_1;
always @(negedge clk)
q40_0<=m40_0;
always @(negedge clk)
q40_1<=m40_1;
always @(negedge clk)
q41_0<=m41_0;
always @(negedge clk)
q41_1<=m41_1;
always @(negedge clk)
q42_0<=m42_0;
always @(negedge clk)
q42_1<=m42_1;
always @(negedge clk)
q43_0<=m43_0;
always @(negedge clk)
q43_1<=m43_1;
always @(negedge clk)
q44_0<=m44_0;
always @(negedge clk)
q44_1<=m44_1;
always @(negedge clk)
q45_0<=m45_0;
always @(negedge clk)
q45_1<=m45_1;
always @(negedge clk)
q46_0<=m46_0;
always @(negedge clk)
q46_1<=m46_1;
always @(negedge clk)
q47_0<=m47_0;
always @(negedge clk)
q47_1<=m47_1;
always @(negedge clk)
q48_0<=m48_0;
always @(negedge clk)
q48_1<=m48_1;
always @(negedge clk)
q49_0<=m49_0;
always @(negedge clk)
q49_1<=m49_1;
always @(negedge clk)
q50_0<=m50_0;
always @(negedge clk)
q50_1<=m50_1;

always @(posedge clk)
m0_0<=h0_0;/*
always @(posedge clk)
m0_1<=h0_1;*/
always @(posedge clk)
m1_0<=h1_0;/*
always @(posedge clk)
m1_1<=h1_1;*/

always @(negedge clk)
q0_0<=m0_0;/*
always @(negedge clk)
q0_1<=m0_1;*/
always @(negedge clk)
q1_0<=m1_0;/*
always @(negedge clk)
q1_1<=m1_1;*/

or     H0000000_0(h0000000_0,h0000000_011,h0000000_012,h0000000_013),
       H0000000_1(h0000000_1,h0000000_111,h0000000_112),
       H0000001_0(h0000001_0,h0000001_011,h0000001_012,h0000001_013),
       H0000001_1(h0000001_1,h0000001_111,h0000001_112),
       H0000010_0(h0000010_0,h0000010_011,h0000010_012,h0000010_013),
       H0000010_1(h0000010_1,h0000010_111,h0000010_112),
       H0000011_0(h0000011_0,h0000011_011,h0000011_012,h0000011_013),
       H0000011_1(h0000011_1,h0000011_111,h0000011_112),
       H0000100_0(h0000100_0,h0000100_011,h0000100_012,h0000100_013),
       H0000100_1(h0000100_1,h0000100_111,h0000100_112),
       H0000101_0(h0000101_0,h0000101_011,h0000101_012,h0000101_013),
       H0000101_1(h0000101_1,h0000101_111,h0000101_112),
       H0000110_0(h0000110_0,h0000110_011,h0000110_012,h0000110_013),
       H0000110_1(h0000110_1,h0000110_111,h0000110_112),
       H0000111_0(h0000111_0,h0000111_011,h0000111_012,h0000111_013),
       H0000111_1(h0000111_1,h0000111_111,h0000111_112),
       H0001000_0(h0001000_0,h0001000_011,h0001000_012,h0001000_013),
       H0001000_1(h0001000_1,h0001000_111,h0001000_112),
       H0001001_0(h0001001_0,h0001001_011,h0001001_012,h0001001_013),
       H0001001_1(h0001001_1,h0001001_111,h0001001_112),
       H0001010_0(h0001010_0,h0001010_011,h0001010_012,h0001010_013),
       H0001010_1(h0001010_1,h0001010_111,h0001010_112),
       H0001011_0(h0001011_0,h0001011_011,h0001011_012,h0001011_013),
       H0001011_1(h0001011_1,h0001011_111,h0001011_112),
       H0001100_0(h0001100_0,h0001100_011,h0001100_012,h0001100_013),
       H0001100_1(h0001100_1,h0001100_111,h0001100_112),
       H0001101_0(h0001101_0,h0001101_011,h0001101_012,h0001101_013),
       H0001101_1(h0001101_1,h0001101_111,h0001101_112),
       H0001110_0(h0001110_0,h0001110_011,h0001110_012,h0001110_013),
       H0001110_1(h0001110_1,h0001110_111,h0001110_112),
       H0001111_0(h0001111_0,h0001111_011,h0001111_012,h0001111_013),
       H0001111_1(h0001111_1,h0001111_111,h0001111_112),
       H0010000_0(h0010000_0,h0010000_011,h0010000_012,h0010000_013),
       H0010000_1(h0010000_1,h0010000_111,h0010000_112),
       H0010001_0(h0010001_0,h0010001_011,h0010001_012,h0010001_013),
       H0010001_1(h0010001_1,h0010001_111,h0010001_112),
       H0010010_0(h0010010_0,h0010010_011,h0010010_012,h0010010_013),
       H0010010_1(h0010010_1,h0010010_111,h0010010_112),
       H0010011_0(h0010011_0,h0010011_011,h0010011_012,h0010011_013),
       H0010011_1(h0010011_1,h0010011_111,h0010011_112),
       H0010100_0(h0010100_0,h0010100_011,h0010100_012,h0010100_013),
       H0010100_1(h0010100_1,h0010100_111,h0010100_112),
       H0010101_0(h0010101_0,h0010101_011,h0010101_012,h0010101_013),
       H0010101_1(h0010101_1,h0010101_111,h0010101_112),
       H0010110_0(h0010110_0,h0010110_011,h0010110_012,h0010110_013),
       H0010110_1(h0010110_1,h0010110_111,h0010110_112),
       H0010111_0(h0010111_0,h0010111_011,h0010111_012,h0010111_013),
       H0010111_1(h0010111_1,h0010111_111,h0010111_112),
       H0011000_0(h0011000_0,h0011000_011,h0011000_012,h0011000_013),
       H0011000_1(h0011000_1,h0011000_111,h0011000_112),
       H0011001_0(h0011001_0,h0011001_011,h0011001_012,h0011001_013),
       H0011001_1(h0011001_1,h0011001_111,h0011001_112),
       H0011010_0(h0011010_0,h0011010_011,h0011010_012,h0011010_013),
       H0011010_1(h0011010_1,h0011010_111,h0011010_112),
       H0011011_0(h0011011_0,h0011011_011,h0011011_012,h0011011_013),
       H0011011_1(h0011011_1,h0011011_111,h0011011_112),
       H0011100_0(h0011100_0,h0011100_011,h0011100_012,h0011100_013),
       H0011100_1(h0011100_1,h0011100_111,h0011100_112),
       H0011101_0(h0011101_0,h0011101_011,h0011101_012,h0011101_013),
       H0011101_1(h0011101_1,h0011101_111,h0011101_112),
       H0011110_0(h0011110_0,h0011110_011,h0011110_012,h0011110_013),
       H0011110_1(h0011110_1,h0011110_111,h0011110_112),
       H0011111_0(h0011111_0,h0011111_011,h0011111_012,h0011111_013),
       H0011111_1(h0011111_1,h0011111_111,h0011111_112),
       H0100000_0(h0100000_0,h0100000_011,h0100000_012,h0100000_013),
       H0100000_1(h0100000_1,h0100000_111,h0100000_112),
       H0100001_0(h0100001_0,h0100001_011,h0100001_012,h0100001_013),
       H0100001_1(h0100001_1,h0100001_111,h0100001_112),
       H0100010_0(h0100010_0,h0100010_011,h0100010_012,h0100010_013),
       H0100010_1(h0100010_1,h0100010_111,h0100010_112),
       H0100011_0(h0100011_0,h0100011_011,h0100011_012,h0100011_013),
       H0100011_1(h0100011_1,h0100011_111,h0100011_112),
       H0100100_0(h0100100_0,h0100100_011,h0100100_012,h0100100_013),
       H0100100_1(h0100100_1,h0100100_111,h0100100_112),
       H0100101_0(h0100101_0,h0100101_011,h0100101_012,h0100101_013),
       H0100101_1(h0100101_1,h0100101_111,h0100101_112),
       H0100110_0(h0100110_0,h0100110_011,h0100110_012,h0100110_013),
       H0100110_1(h0100110_1,h0100110_111,h0100110_112),
       H0100111_0(h0100111_0,h0100111_011,h0100111_012,h0100111_013),
       H0100111_1(h0100111_1,h0100111_111,h0100111_112),
       H0101000_0(h0101000_0,h0101000_011,h0101000_012,h0101000_013),
       H0101000_1(h0101000_1,h0101000_111,h0101000_112),
       H0101001_0(h0101001_0,h0101001_011,h0101001_012,h0101001_013),
       H0101001_1(h0101001_1,h0101001_111,h0101001_112),
       H0101010_0(h0101010_0,h0101010_011,h0101010_012,h0101010_013),
       H0101010_1(h0101010_1,h0101010_111,h0101010_112),
       H0101011_0(h0101011_0,h0101011_011,h0101011_012,h0101011_013),
       H0101011_1(h0101011_1,h0101011_111,h0101011_112),
       H0101100_0(h0101100_0,h0101100_011,h0101100_012,h0101100_013),
       H0101100_1(h0101100_1,h0101100_111,h0101100_112),
       H0101101_0(h0101101_0,h0101101_011,h0101101_012,h0101101_013),
       H0101101_1(h0101101_1,h0101101_111,h0101101_112),
       H0101110_0(h0101110_0,h0101110_011,h0101110_012,h0101110_013),
       H0101110_1(h0101110_1,h0101110_111,h0101110_112),
       H0101111_0(h0101111_0,h0101111_011,h0101111_012,h0101111_013),
       H0101111_1(h0101111_1,h0101111_111,h0101111_112),
       H0110000_0(h0110000_0,h0110000_011,h0110000_012,h0110000_013),
       H0110000_1(h0110000_1,h0110000_111,h0110000_112),
       H0110001_0(h0110001_0,h0110001_011,h0110001_012,h0110001_013),
       H0110001_1(h0110001_1,h0110001_111,h0110001_112),
       H0110010_0(h0110010_0,h0110010_011,h0110010_012,h0110010_013),
       H0110010_1(h0110010_1,h0110010_111,h0110010_112),
       H0110011_0(h0110011_0,h0110011_011,h0110011_012,h0110011_013),
       H0110011_1(h0110011_1,h0110011_111,h0110011_112),
       H0110100_0(h0110100_0,h0110100_011,h0110100_012,h0110100_013),
       H0110100_1(h0110100_1,h0110100_111,h0110100_112),
       H0110101_0(h0110101_0,h0110101_011,h0110101_012,h0110101_013),
       H0110101_1(h0110101_1,h0110101_111,h0110101_112),
       H0110110_0(h0110110_0,h0110110_011,h0110110_012,h0110110_013),
       H0110110_1(h0110110_1,h0110110_111,h0110110_112),
       H0110111_0(h0110111_0,h0110111_011,h0110111_012,h0110111_013),
       H0110111_1(h0110111_1,h0110111_111,h0110111_112),
       H0111000_0(h0111000_0,h0111000_011,h0111000_012,h0111000_013),
       H0111000_1(h0111000_1,h0111000_111,h0111000_112),
       H0111001_0(h0111001_0,h0111001_011,h0111001_012,h0111001_013),
       H0111001_1(h0111001_1,h0111001_111,h0111001_112),
       H0111010_0(h0111010_0,h0111010_011,h0111010_012,h0111010_013),
       H0111010_1(h0111010_1,h0111010_111,h0111010_112),
       H0111011_0(h0111011_0,h0111011_011,h0111011_012,h0111011_013),
       H0111011_1(h0111011_1,h0111011_111,h0111011_112),
       H0111100_0(h0111100_0,h0111100_011,h0111100_012,h0111100_013),
       H0111100_1(h0111100_1,h0111100_111,h0111100_112),
       H0111101_0(h0111101_0,h0111101_011,h0111101_012,h0111101_013),
       H0111101_1(h0111101_1,h0111101_111,h0111101_112),
       H0111110_0(h0111110_0,h0111110_011,h0111110_012,h0111110_013,q11_1),
       H0111110_1(h0111110_1,h0111110_111,h0111110_112,q11_1),
       H0111111_0(h0111111_0,h0111111_011,h0111111_012,h0111111_013,q11_1),
       H0111111_1(h0111111_1,h0111111_111,h0111111_112,q11_1),
       H1000000_0(h1000000_0,h1000000_011,h1000000_012,h1000000_013,q11_1),
       H1000000_1(h1000000_1,h1000000_111,h1000000_112,q11_1),
       H1000001_0(h1000001_0,h1000001_011,h1000001_012,h1000001_013,q11_1),
       H1000001_1(h1000001_1,h1000001_111,h1000001_112,q11_1),
       H1000010_0(h1000010_0,h1000010_011,h1000010_012,h1000010_013),
       H1000010_1(h1000010_1,h1000010_111,h1000010_112),
       H1000011_0(h1000011_0,h1000011_011,h1000011_012,h1000011_013),
       H1000011_1(h1000011_1,h1000011_111,h1000011_112),
       H1000100_0(h1000100_0,h1000100_011,h1000100_012,h1000100_013),
       H1000100_1(h1000100_1,h1000100_111,h1000100_112),
       H1000101_0(h1000101_0,h1000101_011,h1000101_012,h1000101_013),
       H1000101_1(h1000101_1,h1000101_111,h1000101_112),
       H1000110_0(h1000110_0,h1000110_011,h1000110_012,h1000110_013),
       H1000110_1(h1000110_1,h1000110_111,h1000110_112),
       H1000111_0(h1000111_0,h1000111_011,h1000111_012,h1000111_013),
       H1000111_1(h1000111_1,h1000111_111,h1000111_112),
       H1001000_0(h1001000_0,h1001000_011,h1001000_012,h1001000_013),
       H1001000_1(h1001000_1,h1001000_111,h1001000_112),
       H1001001_0(h1001001_0,h1001001_011,h1001001_012,h1001001_013),
       H1001001_1(h1001001_1,h1001001_111,h1001001_112),
       H1001010_0(h1001010_0,h1001010_011,h1001010_012,h1001010_013),
       H1001010_1(h1001010_1,h1001010_111,h1001010_112),
       H1001011_0(h1001011_0,h1001011_011,h1001011_012,h1001011_013),
       H1001011_1(h1001011_1,h1001011_111,h1001011_112),
       H1001100_0(h1001100_0,h1001100_011,h1001100_012,h1001100_013),
       H1001100_1(h1001100_1,h1001100_111,h1001100_112),
       H1001101_0(h1001101_0,h1001101_011,h1001101_012,h1001101_013),
       H1001101_1(h1001101_1,h1001101_111,h1001101_112),
       H1001110_0(h1001110_0,h1001110_011,h1001110_012,h1001110_013),
       H1001110_1(h1001110_1,h1001110_111,h1001110_112),
       H1001111_0(h1001111_0,h1001111_011,h1001111_012,h1001111_013),
       H1001111_1(h1001111_1,h1001111_111,h1001111_112),
       H1010000_0(h1010000_0,h1010000_011,h1010000_012,h1010000_013),
       H1010000_1(h1010000_1,h1010000_111,h1010000_112),
       H1010001_0(h1010001_0,h1010001_011,h1010001_012,h1010001_013),
       H1010001_1(h1010001_1,h1010001_111,h1010001_112),
       H1010010_0(h1010010_0,h1010010_011,h1010010_012,h1010010_013),
       H1010010_1(h1010010_1,h1010010_111,h1010010_112),
       H1010011_0(h1010011_0,h1010011_011,h1010011_012,h1010011_013),
       H1010011_1(h1010011_1,h1010011_111,h1010011_112),
       H1010100_0(h1010100_0,h1010100_011,h1010100_012,h1010100_013),
       H1010100_1(h1010100_1,h1010100_111,h1010100_112),
       H1010101_0(h1010101_0,h1010101_011,h1010101_012,h1010101_013),
       H1010101_1(h1010101_1,h1010101_111,h1010101_112),
       H1010110_0(h1010110_0,h1010110_011,h1010110_012,h1010110_013),
       H1010110_1(h1010110_1,h1010110_111,h1010110_112),
       H1010111_0(h1010111_0,h1010111_011,h1010111_012,h1010111_013),
       H1010111_1(h1010111_1,h1010111_111,h1010111_112),
       H1011000_0(h1011000_0,h1011000_011,h1011000_012,h1011000_013),
       H1011000_1(h1011000_1,h1011000_111,h1011000_112),
       H1011001_0(h1011001_0,h1011001_011,h1011001_012,h1011001_013),
       H1011001_1(h1011001_1,h1011001_111,h1011001_112),
       H1011010_0(h1011010_0,h1011010_011,h1011010_012,h1011010_013),
       H1011010_1(h1011010_1,h1011010_111,h1011010_112),
       H1011011_0(h1011011_0,h1011011_011,h1011011_012,h1011011_013),
       H1011011_1(h1011011_1,h1011011_111,h1011011_112),
       H1011100_0(h1011100_0,h1011100_011,h1011100_012,h1011100_013),
       H1011100_1(h1011100_1,h1011100_111,h1011100_112),
       H1011101_0(h1011101_0,h1011101_011,h1011101_012,h1011101_013),
       H1011101_1(h1011101_1,h1011101_111,h1011101_112),
       H1011110_0(h1011110_0,h1011110_011,h1011110_012,h1011110_013),
       H1011110_1(h1011110_1,h1011110_111,h1011110_112),
       H1011111_0(h1011111_0,h1011111_011,h1011111_012,h1011111_013),
       H1011111_1(h1011111_1,h1011111_111,h1011111_112),
       H1100000_0(h1100000_0,h1100000_011,h1100000_012,h1100000_013),
       H1100000_1(h1100000_1,h1100000_111,h1100000_112),
       H1100001_0(h1100001_0,h1100001_011,h1100001_012,h1100001_013),
       H1100001_1(h1100001_1,h1100001_111,h1100001_112),
       H1100010_0(h1100010_0,h1100010_011,h1100010_012,h1100010_013),
       H1100010_1(h1100010_1,h1100010_111,h1100010_112),
       H1100011_0(h1100011_0,h1100011_011,h1100011_012,h1100011_013),
       H1100011_1(h1100011_1,h1100011_111,h1100011_112),
       H1100100_0(h1100100_0,h1100100_011,h1100100_012,h1100100_013),
       H1100100_1(h1100100_1,h1100100_111,h1100100_112),
       H1100101_0(h1100101_0,h1100101_011,h1100101_012,h1100101_013),
       H1100101_1(h1100101_1,h1100101_111,h1100101_112),
       H1100110_0(h1100110_0,h1100110_011,h1100110_012,h1100110_013),
       H1100110_1(h1100110_1,h1100110_111,h1100110_112),
       H1100111_0(h1100111_0,h1100111_011,h1100111_012,h1100111_013),
       H1100111_1(h1100111_1,h1100111_111,h1100111_112),
       H1101000_0(h1101000_0,h1101000_011,h1101000_012,h1101000_013),
       H1101000_1(h1101000_1,h1101000_111,h1101000_112),
       H1101001_0(h1101001_0,h1101001_011,h1101001_012,h1101001_013),
       H1101001_1(h1101001_1,h1101001_111,h1101001_112),
       H1101010_0(h1101010_0,h1101010_011,h1101010_012,h1101010_013),
       H1101010_1(h1101010_1,h1101010_111,h1101010_112),
       H1101011_0(h1101011_0,h1101011_011,h1101011_012,h1101011_013),
       H1101011_1(h1101011_1,h1101011_111,h1101011_112),
       H1101100_0(h1101100_0,h1101100_011,h1101100_012,h1101100_013),
       H1101100_1(h1101100_1,h1101100_111,h1101100_112),
       H1101101_0(h1101101_0,h1101101_011,h1101101_012,h1101101_013),
       H1101101_1(h1101101_1,h1101101_111,h1101101_112),
       H1101110_0(h1101110_0,h1101110_011,h1101110_012,h1101110_013),
       H1101110_1(h1101110_1,h1101110_111,h1101110_112),
       H1101111_0(h1101111_0,h1101111_011,h1101111_012,h1101111_013),
       H1101111_1(h1101111_1,h1101111_111,h1101111_112),
       H1110000_0(h1110000_0,h1110000_011,h1110000_012,h1110000_013),
       H1110000_1(h1110000_1,h1110000_111,h1110000_112),
       H1110001_0(h1110001_0,h1110001_011,h1110001_012,h1110001_013),
       H1110001_1(h1110001_1,h1110001_111,h1110001_112),
       H1110010_0(h1110010_0,h1110010_011,h1110010_012,h1110010_013),
       H1110010_1(h1110010_1,h1110010_111,h1110010_112),
       H1110011_0(h1110011_0,h1110011_011,h1110011_012,h1110011_013),
       H1110011_1(h1110011_1,h1110011_111,h1110011_112),
       H1110100_0(h1110100_0,h1110100_011,h1110100_012,h1110100_013),
       H1110100_1(h1110100_1,h1110100_111,h1110100_112),
       H1110101_0(h1110101_0,h1110101_011,h1110101_012,h1110101_013),
       H1110101_1(h1110101_1,h1110101_111,h1110101_112),
       H1110110_0(h1110110_0,h1110110_011,h1110110_012,h1110110_013),
       H1110110_1(h1110110_1,h1110110_111,h1110110_112),
       H1110111_0(h1110111_0,h1110111_011,h1110111_012,h1110111_013),
       H1110111_1(h1110111_1,h1110111_111,h1110111_112),
       H1111000_0(h1111000_0,h1111000_011,h1111000_012,h1111000_013),
       H1111000_1(h1111000_1,h1111000_111,h1111000_112),
       H1111001_0(h1111001_0,h1111001_011,h1111001_012,h1111001_013),
       H1111001_1(h1111001_1,h1111001_111,h1111001_112),
       H1111010_0(h1111010_0,h1111010_011,h1111010_012,h1111010_013),
       H1111010_1(h1111010_1,h1111010_111,h1111010_112),
       H1111011_0(h1111011_0,h1111011_011,h1111011_012,h1111011_013),
       H1111011_1(h1111011_1,h1111011_111,h1111011_112),
       H1111100_0(h1111100_0,h1111100_011,h1111100_012,h1111100_013),
       H1111100_1(h1111100_1,h1111100_111,h1111100_112),
       H1111101_0(h1111101_0,h1111101_011,h1111101_012,h1111101_013),
       H1111101_1(h1111101_1,h1111101_111,h1111101_112),
       H1111110_0(h1111110_0,h1111110_011,h1111110_012,h1111110_013),
       H1111110_1(h1111110_1,h1111110_111,h1111110_112),
       H1111111_0(h1111111_0,h1111111_011,h1111111_012,h1111111_013),
       H1111111_1(h1111111_1,h1111111_111,h1111111_112);

and    H0000000_011(h0000000_011,o3190,q0000000_0),
       H0000000_111(h0000000_111,o3190,q0000000_0),
       H0000001_011(h0000001_011,o3190,q0000001_0),
       H0000001_111(h0000001_111,o3190,q0000001_0),
       H0000010_011(h0000010_011,o3190,q0000010_0),
       H0000010_111(h0000010_111,o3190,q0000010_0),
       H0000011_011(h0000011_011,o3190,q0000011_0),
       H0000011_111(h0000011_111,o3190,q0000011_0),
       H0000100_011(h0000100_011,o3190,q0000100_0),
       H0000100_111(h0000100_111,o3190,q0000100_0),
       H0000101_011(h0000101_011,o3190,q0000101_0),
       H0000101_111(h0000101_111,o3190,q0000101_0),
       H0000110_011(h0000110_011,o3190,q0000110_0),
       H0000110_111(h0000110_111,o3190,q0000110_0),
       H0000111_011(h0000111_011,o3190,q0000111_0),
       H0000111_111(h0000111_111,o3190,q0000111_0),
       H0001000_011(h0001000_011,o3190,q0001000_0),
       H0001000_111(h0001000_111,o3190,q0001000_0),
       H0001001_011(h0001001_011,o3190,q0001001_0),
       H0001001_111(h0001001_111,o3190,q0001001_0),
       H0001010_011(h0001010_011,o3190,q0001010_0),
       H0001010_111(h0001010_111,o3190,q0001010_0),
       H0001011_011(h0001011_011,o3190,q0001011_0),
       H0001011_111(h0001011_111,o3190,q0001011_0),
       H0001100_011(h0001100_011,o3190,q0001100_0),
       H0001100_111(h0001100_111,o3190,q0001100_0),
       H0001101_011(h0001101_011,o3190,q0001101_0),
       H0001101_111(h0001101_111,o3190,q0001101_0),
       H0001110_011(h0001110_011,o3190,q0001110_0),
       H0001110_111(h0001110_111,o3190,q0001110_0),
       H0001111_011(h0001111_011,o3190,q0001111_0),
       H0001111_111(h0001111_111,o3190,q0001111_0),
       H0010000_011(h0010000_011,o3190,q0010000_0),
       H0010000_111(h0010000_111,o3190,q0010000_0),
       H0010001_011(h0010001_011,o3190,q0010001_0),
       H0010001_111(h0010001_111,o3190,q0010001_0),
       H0010010_011(h0010010_011,o3190,q0010010_0),
       H0010010_111(h0010010_111,o3190,q0010010_0),
       H0010011_011(h0010011_011,o3190,q0010011_0),
       H0010011_111(h0010011_111,o3190,q0010011_0),
       H0010100_011(h0010100_011,o3190,q0010100_0),
       H0010100_111(h0010100_111,o3190,q0010100_0),
       H0010101_011(h0010101_011,o3190,q0010101_0),
       H0010101_111(h0010101_111,o3190,q0010101_0),
       H0010110_011(h0010110_011,o3190,q0010110_0),
       H0010110_111(h0010110_111,o3190,q0010110_0),
       H0010111_011(h0010111_011,o3190,q0010111_0),
       H0010111_111(h0010111_111,o3190,q0010111_0),
       H0011000_011(h0011000_011,o3190,q0011000_0),
       H0011000_111(h0011000_111,o3190,q0011000_0),
       H0011001_011(h0011001_011,o3190,q0011001_0),
       H0011001_111(h0011001_111,o3190,q0011001_0),
       H0011010_011(h0011010_011,o3190,q0011010_0),
       H0011010_111(h0011010_111,o3190,q0011010_0),
       H0011011_011(h0011011_011,o3190,q0011011_0),
       H0011011_111(h0011011_111,o3190,q0011011_0),
       H0011100_011(h0011100_011,o3190,q0011100_0),
       H0011100_111(h0011100_111,o3190,q0011100_0),
       H0011101_011(h0011101_011,o3190,q0011101_0),
       H0011101_111(h0011101_111,o3190,q0011101_0),
       H0011110_011(h0011110_011,o3190,q0011110_0),
       H0011110_111(h0011110_111,o3190,q0011110_0),
       H0011111_011(h0011111_011,o3190,q0011111_0),
       H0011111_111(h0011111_111,o3190,q0011111_0),
       H0100000_011(h0100000_011,o3190,q0100000_0),
       H0100000_111(h0100000_111,o3190,q0100000_0),
       H0100001_011(h0100001_011,o3190,q0100001_0),
       H0100001_111(h0100001_111,o3190,q0100001_0),
       H0100010_011(h0100010_011,o3190,q0100010_0),
       H0100010_111(h0100010_111,o3190,q0100010_0),
       H0100011_011(h0100011_011,o3190,q0100011_0),
       H0100011_111(h0100011_111,o3190,q0100011_0),
       H0100100_011(h0100100_011,o3190,q0100100_0),
       H0100100_111(h0100100_111,o3190,q0100100_0),
       H0100101_011(h0100101_011,o3190,q0100101_0),
       H0100101_111(h0100101_111,o3190,q0100101_0),
       H0100110_011(h0100110_011,o3190,q0100110_0),
       H0100110_111(h0100110_111,o3190,q0100110_0),
       H0100111_011(h0100111_011,o3190,q0100111_0),
       H0100111_111(h0100111_111,o3190,q0100111_0),
       H0101000_011(h0101000_011,o3190,q0101000_0),
       H0101000_111(h0101000_111,o3190,q0101000_0),
       H0101001_011(h0101001_011,o3190,q0101001_0),
       H0101001_111(h0101001_111,o3190,q0101001_0),
       H0101010_011(h0101010_011,o3190,q0101010_0),
       H0101010_111(h0101010_111,o3190,q0101010_0),
       H0101011_011(h0101011_011,o3190,q0101011_0),
       H0101011_111(h0101011_111,o3190,q0101011_0),
       H0101100_011(h0101100_011,o3190,q0101100_0),
       H0101100_111(h0101100_111,o3190,q0101100_0),
       H0101101_011(h0101101_011,o3190,q0101101_0),
       H0101101_111(h0101101_111,o3190,q0101101_0),
       H0101110_011(h0101110_011,o3190,q0101110_0),
       H0101110_111(h0101110_111,o3190,q0101110_0),
       H0101111_011(h0101111_011,o3190,q0101111_0),
       H0101111_111(h0101111_111,o3190,q0101111_0),
       H0110000_011(h0110000_011,o3190,q0110000_0),
       H0110000_111(h0110000_111,o3190,q0110000_0),
       H0110001_011(h0110001_011,o3190,q0110001_0),
       H0110001_111(h0110001_111,o3190,q0110001_0),
       H0110010_011(h0110010_011,o3190,q0110010_0),
       H0110010_111(h0110010_111,o3190,q0110010_0),
       H0110011_011(h0110011_011,o3190,q0110011_0),
       H0110011_111(h0110011_111,o3190,q0110011_0),
       H0110100_011(h0110100_011,o3190,q0110100_0),
       H0110100_111(h0110100_111,o3190,q0110100_0),
       H0110101_011(h0110101_011,o3190,q0110101_0),
       H0110101_111(h0110101_111,o3190,q0110101_0),
       H0110110_011(h0110110_011,o3190,q0110110_0),
       H0110110_111(h0110110_111,o3190,q0110110_0),
       H0110111_011(h0110111_011,o3190,q0110111_0),
       H0110111_111(h0110111_111,o3190,q0110111_0),
       H0111000_011(h0111000_011,o3190,q0111000_0),
       H0111000_111(h0111000_111,o3190,q0111000_0),
       H0111001_011(h0111001_011,o3190,q0111001_0),
       H0111001_111(h0111001_111,o3190,q0111001_0),
       H0111010_011(h0111010_011,o3190,q0111010_0),
       H0111010_111(h0111010_111,o3190,q0111010_0),
       H0111011_011(h0111011_011,o3190,q0111011_0),
       H0111011_111(h0111011_111,o3190,q0111011_0),
       H0111100_011(h0111100_011,o3190,q0111100_0),
       H0111100_111(h0111100_111,o3190,q0111100_0),
       H0111101_011(h0111101_011,o3190,q0111101_0),
       H0111101_111(h0111101_111,o3190,q0111101_0),
       H0111110_011(h0111110_011,o3190,q0111110_0),
       H0111110_111(h0111110_111,o3190,q0111110_0),
       H0111111_011(h0111111_011,o3190,q0111111_0),
       H0111111_111(h0111111_111,o3190,q0111111_0),
       H1000000_011(h1000000_011,o3190,q1000000_0),
       H1000000_111(h1000000_111,o3190,q1000000_0),
       H1000001_011(h1000001_011,o3190,q1000001_0),
       H1000001_111(h1000001_111,o3190,q1000001_0),
       H1000010_011(h1000010_011,o3190,q1000010_0),
       H1000010_111(h1000010_111,o3190,q1000010_0),
       H1000011_011(h1000011_011,o3190,q1000011_0),
       H1000011_111(h1000011_111,o3190,q1000011_0),
       H1000100_011(h1000100_011,o3190,q1000100_0),
       H1000100_111(h1000100_111,o3190,q1000100_0),
       H1000101_011(h1000101_011,o3190,q1000101_0),
       H1000101_111(h1000101_111,o3190,q1000101_0),
       H1000110_011(h1000110_011,o3190,q1000110_0),
       H1000110_111(h1000110_111,o3190,q1000110_0),
       H1000111_011(h1000111_011,o3190,q1000111_0),
       H1000111_111(h1000111_111,o3190,q1000111_0),
       H1001000_011(h1001000_011,o3190,q1001000_0),
       H1001000_111(h1001000_111,o3190,q1001000_0),
       H1001001_011(h1001001_011,o3190,q1001001_0),
       H1001001_111(h1001001_111,o3190,q1001001_0),
       H1001010_011(h1001010_011,o3190,q1001010_0),
       H1001010_111(h1001010_111,o3190,q1001010_0),
       H1001011_011(h1001011_011,o3190,q1001011_0),
       H1001011_111(h1001011_111,o3190,q1001011_0),
       H1001100_011(h1001100_011,o3190,q1001100_0),
       H1001100_111(h1001100_111,o3190,q1001100_0),
       H1001101_011(h1001101_011,o3190,q1001101_0),
       H1001101_111(h1001101_111,o3190,q1001101_0),
       H1001110_011(h1001110_011,o3190,q1001110_0),
       H1001110_111(h1001110_111,o3190,q1001110_0),
       H1001111_011(h1001111_011,o3190,q1001111_0),
       H1001111_111(h1001111_111,o3190,q1001111_0),
       H1010000_011(h1010000_011,o3190,q1010000_0),
       H1010000_111(h1010000_111,o3190,q1010000_0),
       H1010001_011(h1010001_011,o3190,q1010001_0),
       H1010001_111(h1010001_111,o3190,q1010001_0),
       H1010010_011(h1010010_011,o3190,q1010010_0),
       H1010010_111(h1010010_111,o3190,q1010010_0),
       H1010011_011(h1010011_011,o3190,q1010011_0),
       H1010011_111(h1010011_111,o3190,q1010011_0),
       H1010100_011(h1010100_011,o3190,q1010100_0),
       H1010100_111(h1010100_111,o3190,q1010100_0),
       H1010101_011(h1010101_011,o3190,q1010101_0),
       H1010101_111(h1010101_111,o3190,q1010101_0),
       H1010110_011(h1010110_011,o3190,q1010110_0),
       H1010110_111(h1010110_111,o3190,q1010110_0),
       H1010111_011(h1010111_011,o3190,q1010111_0),
       H1010111_111(h1010111_111,o3190,q1010111_0),
       H1011000_011(h1011000_011,o3190,q1011000_0),
       H1011000_111(h1011000_111,o3190,q1011000_0),
       H1011001_011(h1011001_011,o3190,q1011001_0),
       H1011001_111(h1011001_111,o3190,q1011001_0),
       H1011010_011(h1011010_011,o3190,q1011010_0),
       H1011010_111(h1011010_111,o3190,q1011010_0),
       H1011011_011(h1011011_011,o3190,q1011011_0),
       H1011011_111(h1011011_111,o3190,q1011011_0),
       H1011100_011(h1011100_011,o3190,q1011100_0),
       H1011100_111(h1011100_111,o3190,q1011100_0),
       H1011101_011(h1011101_011,o3190,q1011101_0),
       H1011101_111(h1011101_111,o3190,q1011101_0),
       H1011110_011(h1011110_011,o3190,q1011110_0),
       H1011110_111(h1011110_111,o3190,q1011110_0),
       H1011111_011(h1011111_011,o3190,q1011111_0),
       H1011111_111(h1011111_111,o3190,q1011111_0),
       H1100000_011(h1100000_011,o3190,q1100000_0),
       H1100000_111(h1100000_111,o3190,q1100000_0),
       H1100001_011(h1100001_011,o3190,q1100001_0),
       H1100001_111(h1100001_111,o3190,q1100001_0),
       H1100010_011(h1100010_011,o3190,q1100010_0),
       H1100010_111(h1100010_111,o3190,q1100010_0),
       H1100011_011(h1100011_011,o3190,q1100011_0),
       H1100011_111(h1100011_111,o3190,q1100011_0),
       H1100100_011(h1100100_011,o3190,q1100100_0),
       H1100100_111(h1100100_111,o3190,q1100100_0),
       H1100101_011(h1100101_011,o3190,q1100101_0),
       H1100101_111(h1100101_111,o3190,q1100101_0),
       H1100110_011(h1100110_011,o3190,q1100110_0),
       H1100110_111(h1100110_111,o3190,q1100110_0),
       H1100111_011(h1100111_011,o3190,q1100111_0),
       H1100111_111(h1100111_111,o3190,q1100111_0),
       H1101000_011(h1101000_011,o3190,q1101000_0),
       H1101000_111(h1101000_111,o3190,q1101000_0),
       H1101001_011(h1101001_011,o3190,q1101001_0),
       H1101001_111(h1101001_111,o3190,q1101001_0),
       H1101010_011(h1101010_011,o3190,q1101010_0),
       H1101010_111(h1101010_111,o3190,q1101010_0),
       H1101011_011(h1101011_011,o3190,q1101011_0),
       H1101011_111(h1101011_111,o3190,q1101011_0),
       H1101100_011(h1101100_011,o3190,q1101100_0),
       H1101100_111(h1101100_111,o3190,q1101100_0),
       H1101101_011(h1101101_011,o3190,q1101101_0),
       H1101101_111(h1101101_111,o3190,q1101101_0),
       H1101110_011(h1101110_011,o3190,q1101110_0),
       H1101110_111(h1101110_111,o3190,q1101110_0),
       H1101111_011(h1101111_011,o3190,q1101111_0),
       H1101111_111(h1101111_111,o3190,q1101111_0),
       H1110000_011(h1110000_011,o3190,q1110000_0),
       H1110000_111(h1110000_111,o3190,q1110000_0),
       H1110001_011(h1110001_011,o3190,q1110001_0),
       H1110001_111(h1110001_111,o3190,q1110001_0),
       H1110010_011(h1110010_011,o3190,q1110010_0),
       H1110010_111(h1110010_111,o3190,q1110010_0),
       H1110011_011(h1110011_011,o3190,q1110011_0),
       H1110011_111(h1110011_111,o3190,q1110011_0),
       H1110100_011(h1110100_011,o3190,q1110100_0),
       H1110100_111(h1110100_111,o3190,q1110100_0),
       H1110101_011(h1110101_011,o3190,q1110101_0),
       H1110101_111(h1110101_111,o3190,q1110101_0),
       H1110110_011(h1110110_011,o3190,q1110110_0),
       H1110110_111(h1110110_111,o3190,q1110110_0),
       H1110111_011(h1110111_011,o3190,q1110111_0),
       H1110111_111(h1110111_111,o3190,q1110111_0),
       H1111000_011(h1111000_011,o3190,q1111000_0),
       H1111000_111(h1111000_111,o3190,q1111000_0),
       H1111001_011(h1111001_011,o3190,q1111001_0),
       H1111001_111(h1111001_111,o3190,q1111001_0),
       H1111010_011(h1111010_011,o3190,q1111010_0),
       H1111010_111(h1111010_111,o3190,q1111010_0),
       H1111011_011(h1111011_011,o3190,q1111011_0),
       H1111011_111(h1111011_111,o3190,q1111011_0),
       H1111100_011(h1111100_011,o3190,q1111100_0),
       H1111100_111(h1111100_111,o3190,q1111100_0),
       H1111101_011(h1111101_011,o3190,q1111101_0),
       H1111101_111(h1111101_111,o3190,q1111101_0),
       H1111110_011(h1111110_011,o3190,q1111110_0),
       H1111110_111(h1111110_111,o3190,q1111110_0),
       H1111111_011(h1111111_011,o3190,q1111111_0),
       H1111111_111(h1111111_111,o3190,q1111111_0),
       H0000000_012(h0000000_012,n3190,q0_0,dbv0),
       H0000000_112(h0000000_112,n3190,q0000000_1),
       H0000001_012(h0000001_012,n3190,q0_0,q0000000_1),
       H0000001_112(h0000001_112,n3190,q0000001_1),
       H0000010_012(h0000010_012,n3190,q0_0,q0000001_1),
       H0000010_112(h0000010_112,n3190,q0000010_1),
       H0000011_012(h0000011_012,n3190,q0_0,q0000010_1),
       H0000011_112(h0000011_112,n3190,q0000011_1),
       H0000100_012(h0000100_012,n3190,q0_0,q0000011_1),
       H0000100_112(h0000100_112,n3190,q0000100_1),
       H0000101_012(h0000101_012,n3190,q0_0,q0000100_1),
       H0000101_112(h0000101_112,n3190,q0000101_1),
       H0000110_012(h0000110_012,n3190,q0_0,q0000101_1),
       H0000110_112(h0000110_112,n3190,q0000110_1),
       H0000111_012(h0000111_012,n3190,q0_0,q0000110_1),
       H0000111_112(h0000111_112,n3190,q0000111_1),
       H0001000_012(h0001000_012,n3190,q0_0,q0000111_1),
       H0001000_112(h0001000_112,n3190,q0001000_1),
       H0001001_012(h0001001_012,n3190,q0_0,q0001000_1),
       H0001001_112(h0001001_112,n3190,q0001001_1),
       H0001010_012(h0001010_012,n3190,q0_0,q0001001_1),
       H0001010_112(h0001010_112,n3190,q0001010_1),
       H0001011_012(h0001011_012,n3190,q0_0,q0001010_1),
       H0001011_112(h0001011_112,n3190,q0001011_1),
       H0001100_012(h0001100_012,n3190,q0_0,q0001011_1),
       H0001100_112(h0001100_112,n3190,q0001100_1),
       H0001101_012(h0001101_012,n3190,q0_0,q0001100_1),
       H0001101_112(h0001101_112,n3190,q0001101_1),
       H0001110_012(h0001110_012,n3190,q0_0,q0001101_1),
       H0001110_112(h0001110_112,n3190,q0001110_1),
       H0001111_012(h0001111_012,n3190,q0_0,q0001110_1),
       H0001111_112(h0001111_112,n3190,q0001111_1),
       H0010000_012(h0010000_012,n3190,q0_0,q0001111_1),
       H0010000_112(h0010000_112,n3190,q0010000_1),
       H0010001_012(h0010001_012,n3190,q0_0,q0010000_1),
       H0010001_112(h0010001_112,n3190,q0010001_1),
       H0010010_012(h0010010_012,n3190,q0_0,q0010001_1),
       H0010010_112(h0010010_112,n3190,q0010010_1),
       H0010011_012(h0010011_012,n3190,q0_0,q0010010_1),
       H0010011_112(h0010011_112,n3190,q0010011_1),
       H0010100_012(h0010100_012,n3190,q0_0,q0010011_1),
       H0010100_112(h0010100_112,n3190,q0010100_1),
       H0010101_012(h0010101_012,n3190,q0_0,q0010100_1),
       H0010101_112(h0010101_112,n3190,q0010101_1),
       H0010110_012(h0010110_012,n3190,q0_0,q0010101_1),
       H0010110_112(h0010110_112,n3190,q0010110_1),
       H0010111_012(h0010111_012,n3190,q0_0,q0010110_1),
       H0010111_112(h0010111_112,n3190,q0010111_1),
       H0011000_012(h0011000_012,n3190,q0_0,q0010111_1),
       H0011000_112(h0011000_112,n3190,q0011000_1),
       H0011001_012(h0011001_012,n3190,q0_0,q0011000_1),
       H0011001_112(h0011001_112,n3190,q0011001_1),
       H0011010_012(h0011010_012,n3190,q0_0,q0011001_1),
       H0011010_112(h0011010_112,n3190,q0011010_1),
       H0011011_012(h0011011_012,n3190,q0_0,q0011010_1),
       H0011011_112(h0011011_112,n3190,q0011011_1),
       H0011100_012(h0011100_012,n3190,q0_0,q0011011_1),
       H0011100_112(h0011100_112,n3190,q0011100_1),
       H0011101_012(h0011101_012,n3190,q0_0,q0011100_1),
       H0011101_112(h0011101_112,n3190,q0011101_1),
       H0011110_012(h0011110_012,n3190,q0_0,q0011101_1),
       H0011110_112(h0011110_112,n3190,q0011110_1),
       H0011111_012(h0011111_012,n3190,q0_0,q0011110_1),
       H0011111_112(h0011111_112,n3190,q0011111_1),
       H0100000_012(h0100000_012,n3190,q0_0,q0011111_1),
       H0100000_112(h0100000_112,n3190,q0100000_1),
       H0100001_012(h0100001_012,n3190,q0_0,q0100000_1),
       H0100001_112(h0100001_112,n3190,q0100001_1),
       H0100010_012(h0100010_012,n3190,q0_0,q0100001_1),
       H0100010_112(h0100010_112,n3190,q0100010_1),
       H0100011_012(h0100011_012,n3190,q0_0,q0100010_1),
       H0100011_112(h0100011_112,n3190,q0100011_1),
       H0100100_012(h0100100_012,n3190,q0_0,q0100011_1),
       H0100100_112(h0100100_112,n3190,q0100100_1),
       H0100101_012(h0100101_012,n3190,q0_0,q0100100_1),
       H0100101_112(h0100101_112,n3190,q0100101_1),
       H0100110_012(h0100110_012,n3190,q0_0,q0100101_1),
       H0100110_112(h0100110_112,n3190,q0100110_1),
       H0100111_012(h0100111_012,n3190,q0_0,q0100110_1),
       H0100111_112(h0100111_112,n3190,q0100111_1),
       H0101000_012(h0101000_012,n3190,q0_0,q0100111_1),
       H0101000_112(h0101000_112,n3190,q0101000_1),
       H0101001_012(h0101001_012,n3190,q0_0,q0101000_1),
       H0101001_112(h0101001_112,n3190,q0101001_1),
       H0101010_012(h0101010_012,n3190,q0_0,q0101001_1),
       H0101010_112(h0101010_112,n3190,q0101010_1),
       H0101011_012(h0101011_012,n3190,q0_0,q0101010_1),
       H0101011_112(h0101011_112,n3190,q0101011_1),
       H0101100_012(h0101100_012,n3190,q0_0,q0101011_1),
       H0101100_112(h0101100_112,n3190,q0101100_1),
       H0101101_012(h0101101_012,n3190,q0_0,q0101100_1),
       H0101101_112(h0101101_112,n3190,q0101101_1),
       H0101110_012(h0101110_012,n3190,q0_0,q0101101_1),
       H0101110_112(h0101110_112,n3190,q0101110_1),
       H0101111_012(h0101111_012,n3190,q0_0,q0101110_1),
       H0101111_112(h0101111_112,n3190,q0101111_1),
       H0110000_012(h0110000_012,n3190,q0_0,q0101111_1),
       H0110000_112(h0110000_112,n3190,q0110000_1),
       H0110001_012(h0110001_012,n3190,q0_0,q0110000_1),
       H0110001_112(h0110001_112,n3190,q0110001_1),
       H0110010_012(h0110010_012,n3190,q0_0,q0110001_1),
       H0110010_112(h0110010_112,n3190,q0110010_1),
       H0110011_012(h0110011_012,n3190,q0_0,q0110010_1),
       H0110011_112(h0110011_112,n3190,q0110011_1),
       H0110100_012(h0110100_012,n3190,q0_0,q0110011_1),
       H0110100_112(h0110100_112,n3190,q0110100_1),
       H0110101_012(h0110101_012,n3190,q0_0,q0110100_1),
       H0110101_112(h0110101_112,n3190,q0110101_1),
       H0110110_012(h0110110_012,n3190,q0_0,q0110101_1),
       H0110110_112(h0110110_112,n3190,q0110110_1),
       H0110111_012(h0110111_012,n3190,q0_0,q0110110_1),
       H0110111_112(h0110111_112,n3190,q0110111_1),
       H0111000_012(h0111000_012,n3190,q0_0,q0110111_1),
       H0111000_112(h0111000_112,n3190,q0111000_1),
       H0111001_012(h0111001_012,n3190,q0_0,q0111000_1),
       H0111001_112(h0111001_112,n3190,q0111001_1),
       H0111010_012(h0111010_012,n3190,q0_0,q0111001_1),
       H0111010_112(h0111010_112,n3190,q0111010_1),
       H0111011_012(h0111011_012,n3190,q0_0,q0111010_1),
       H0111011_112(h0111011_112,n3190,q0111011_1),
       H0111100_012(h0111100_012,n3190,q0_0,q0111011_1),
       H0111100_112(h0111100_112,n3190,q0111100_1),
       H0111101_012(h0111101_012,n3190,q0_0,q0111100_1),
       H0111101_112(h0111101_112,n3190,q0111101_1),
       H0111110_012(h0111110_012,n3190,q0_0,q0111101_1),
       H0111110_112(h0111110_112,n3190,q0111110_1),
       H0111111_012(h0111111_012,n3190,q0_0,q0111110_1),
       H0111111_112(h0111111_112,n3190,q0111111_1),
       H1000000_012(h1000000_012,n3190,q0_0,q0111111_1),
       H1000000_112(h1000000_112,n3190,q1000000_1),
       H1000001_012(h1000001_012,n3190,q0_0,q1000000_1),
       H1000001_112(h1000001_112,n3190,q1000001_1),
       H1000010_012(h1000010_012,n3190,q0_0,q1000001_1),
       H1000010_112(h1000010_112,n3190,q1000010_1),
       H1000011_012(h1000011_012,n3190,q0_0,q1000010_1),
       H1000011_112(h1000011_112,n3190,q1000011_1),
       H1000100_012(h1000100_012,n3190,q0_0,q1000011_1),
       H1000100_112(h1000100_112,n3190,q1000100_1),
       H1000101_012(h1000101_012,n3190,q0_0,q1000100_1),
       H1000101_112(h1000101_112,n3190,q1000101_1),
       H1000110_012(h1000110_012,n3190,q0_0,q1000101_1),
       H1000110_112(h1000110_112,n3190,q1000110_1),
       H1000111_012(h1000111_012,n3190,q0_0,q1000110_1),
       H1000111_112(h1000111_112,n3190,q1000111_1),
       H1001000_012(h1001000_012,n3190,q0_0,q1000111_1),
       H1001000_112(h1001000_112,n3190,q1001000_1),
       H1001001_012(h1001001_012,n3190,q0_0,q1001000_1),
       H1001001_112(h1001001_112,n3190,q1001001_1),
       H1001010_012(h1001010_012,n3190,q0_0,q1001001_1),
       H1001010_112(h1001010_112,n3190,q1001010_1),
       H1001011_012(h1001011_012,n3190,q0_0,q1001010_1),
       H1001011_112(h1001011_112,n3190,q1001011_1),
       H1001100_012(h1001100_012,n3190,q0_0,q1001011_1),
       H1001100_112(h1001100_112,n3190,q1001100_1),
       H1001101_012(h1001101_012,n3190,q0_0,q1001100_1),
       H1001101_112(h1001101_112,n3190,q1001101_1),
       H1001110_012(h1001110_012,n3190,q0_0,q1001101_1),
       H1001110_112(h1001110_112,n3190,q1001110_1),
       H1001111_012(h1001111_012,n3190,q0_0,q1001110_1),
       H1001111_112(h1001111_112,n3190,q1001111_1),
       H1010000_012(h1010000_012,n3190,q0_0,q1001111_1),
       H1010000_112(h1010000_112,n3190,q1010000_1),
       H1010001_012(h1010001_012,n3190,q0_0,q1010000_1),
       H1010001_112(h1010001_112,n3190,q1010001_1),
       H1010010_012(h1010010_012,n3190,q0_0,q1010001_1),
       H1010010_112(h1010010_112,n3190,q1010010_1),
       H1010011_012(h1010011_012,n3190,q0_0,q1010010_1),
       H1010011_112(h1010011_112,n3190,q1010011_1),
       H1010100_012(h1010100_012,n3190,q0_0,q1010011_1),
       H1010100_112(h1010100_112,n3190,q1010100_1),
       H1010101_012(h1010101_012,n3190,q0_0,q1010100_1),
       H1010101_112(h1010101_112,n3190,q1010101_1),
       H1010110_012(h1010110_012,n3190,q0_0,q1010101_1),
       H1010110_112(h1010110_112,n3190,q1010110_1),
       H1010111_012(h1010111_012,n3190,q0_0,q1010110_1),
       H1010111_112(h1010111_112,n3190,q1010111_1),
       H1011000_012(h1011000_012,n3190,q0_0,q1010111_1),
       H1011000_112(h1011000_112,n3190,q1011000_1),
       H1011001_012(h1011001_012,n3190,q0_0,q1011000_1),
       H1011001_112(h1011001_112,n3190,q1011001_1),
       H1011010_012(h1011010_012,n3190,q0_0,q1011001_1),
       H1011010_112(h1011010_112,n3190,q1011010_1),
       H1011011_012(h1011011_012,n3190,q0_0,q1011010_1),
       H1011011_112(h1011011_112,n3190,q1011011_1),
       H1011100_012(h1011100_012,n3190,q0_0,q1011011_1),
       H1011100_112(h1011100_112,n3190,q1011100_1),
       H1011101_012(h1011101_012,n3190,q0_0,q1011100_1),
       H1011101_112(h1011101_112,n3190,q1011101_1),
       H1011110_012(h1011110_012,n3190,q0_0,q1011101_1),
       H1011110_112(h1011110_112,n3190,q1011110_1),
       H1011111_012(h1011111_012,n3190,q0_0,q1011110_1),
       H1011111_112(h1011111_112,n3190,q1011111_1),
       H1100000_012(h1100000_012,n3190,q0_0,q1011111_1),
       H1100000_112(h1100000_112,n3190,q1100000_1),
       H1100001_012(h1100001_012,n3190,q0_0,q1100000_1),
       H1100001_112(h1100001_112,n3190,q1100001_1),
       H1100010_012(h1100010_012,n3190,q0_0,q1100001_1),
       H1100010_112(h1100010_112,n3190,q1100010_1),
       H1100011_012(h1100011_012,n3190,q0_0,q1100010_1),
       H1100011_112(h1100011_112,n3190,q1100011_1),
       H1100100_012(h1100100_012,n3190,q0_0,q1100011_1),
       H1100100_112(h1100100_112,n3190,q1100100_1),
       H1100101_012(h1100101_012,n3190,q0_0,q1100100_1),
       H1100101_112(h1100101_112,n3190,q1100101_1),
       H1100110_012(h1100110_012,n3190,q0_0,q1100101_1),
       H1100110_112(h1100110_112,n3190,q1100110_1),
       H1100111_012(h1100111_012,n3190,q0_0,q1100110_1),
       H1100111_112(h1100111_112,n3190,q1100111_1),
       H1101000_012(h1101000_012,n3190,q0_0,q1100111_1),
       H1101000_112(h1101000_112,n3190,q1101000_1),
       H1101001_012(h1101001_012,n3190,q0_0,q1101000_1),
       H1101001_112(h1101001_112,n3190,q1101001_1),
       H1101010_012(h1101010_012,n3190,q0_0,q1101001_1),
       H1101010_112(h1101010_112,n3190,q1101010_1),
       H1101011_012(h1101011_012,n3190,q0_0,q1101010_1),
       H1101011_112(h1101011_112,n3190,q1101011_1),
       H1101100_012(h1101100_012,n3190,q0_0,q1101011_1),
       H1101100_112(h1101100_112,n3190,q1101100_1),
       H1101101_012(h1101101_012,n3190,q0_0,q1101100_1),
       H1101101_112(h1101101_112,n3190,q1101101_1),
       H1101110_012(h1101110_012,n3190,q0_0,q1101101_1),
       H1101110_112(h1101110_112,n3190,q1101110_1),
       H1101111_012(h1101111_012,n3190,q0_0,q1101110_1),
       H1101111_112(h1101111_112,n3190,q1101111_1),
       H1110000_012(h1110000_012,n3190,q0_0,q1101111_1),
       H1110000_112(h1110000_112,n3190,q1110000_1),
       H1110001_012(h1110001_012,n3190,q0_0,q1110000_1),
       H1110001_112(h1110001_112,n3190,q1110001_1),
       H1110010_012(h1110010_012,n3190,q0_0,q1110001_1),
       H1110010_112(h1110010_112,n3190,q1110010_1),
       H1110011_012(h1110011_012,n3190,q0_0,q1110010_1),
       H1110011_112(h1110011_112,n3190,q1110011_1),
       H1110100_012(h1110100_012,n3190,q0_0,q1110011_1),
       H1110100_112(h1110100_112,n3190,q1110100_1),
       H1110101_012(h1110101_012,n3190,q0_0,q1110100_1),
       H1110101_112(h1110101_112,n3190,q1110101_1),
       H1110110_012(h1110110_012,n3190,q0_0,q1110101_1),
       H1110110_112(h1110110_112,n3190,q1110110_1),
       H1110111_012(h1110111_012,n3190,q0_0,q1110110_1),
       H1110111_112(h1110111_112,n3190,q1110111_1),
       H1111000_012(h1111000_012,n3190,q0_0,q1110111_1),
       H1111000_112(h1111000_112,n3190,q1111000_1),
       H1111001_012(h1111001_012,n3190,q0_0,q1111000_1),
       H1111001_112(h1111001_112,n3190,q1111001_1),
       H1111010_012(h1111010_012,n3190,q0_0,q1111001_1),
       H1111010_112(h1111010_112,n3190,q1111010_1),
       H1111011_012(h1111011_012,n3190,q0_0,q1111010_1),
       H1111011_112(h1111011_112,n3190,q1111011_1),
       H1111100_012(h1111100_012,n3190,q0_0,q1111011_1),
       H1111100_112(h1111100_112,n3190,q1111100_1),
       H1111101_012(h1111101_012,n3190,q0_0,q1111100_1),
       H1111101_112(h1111101_112,n3190,q1111101_1),
       H1111110_012(h1111110_012,n3190,q0_0,q1111101_1),
       H1111110_112(h1111110_112,n3190,q1111110_1),
       H1111111_012(h1111111_012,n3190,q0_0,q1111110_1),
       H1111111_112(h1111111_112,n3190,q1111111_1),
       H0000000_013(h0000000_013,n3190,n0_0,q0000001_1),
       H0000001_013(h0000001_013,n3190,n0_0,q0000010_1),
       H0000010_013(h0000010_013,n3190,n0_0,q0000011_1),
       H0000011_013(h0000011_013,n3190,n0_0,q0000100_1),
       H0000100_013(h0000100_013,n3190,n0_0,q0000101_1),
       H0000101_013(h0000101_013,n3190,n0_0,q0000110_1),
       H0000110_013(h0000110_013,n3190,n0_0,q0000111_1),
       H0000111_013(h0000111_013,n3190,n0_0,q0001000_1),
       H0001000_013(h0001000_013,n3190,n0_0,q0001001_1),
       H0001001_013(h0001001_013,n3190,n0_0,q0001010_1),
       H0001010_013(h0001010_013,n3190,n0_0,q0001011_1),
       H0001011_013(h0001011_013,n3190,n0_0,q0001100_1),
       H0001100_013(h0001100_013,n3190,n0_0,q0001101_1),
       H0001101_013(h0001101_013,n3190,n0_0,q0001110_1),
       H0001110_013(h0001110_013,n3190,n0_0,q0001111_1),
       H0001111_013(h0001111_013,n3190,n0_0,q0010000_1),
       H0010000_013(h0010000_013,n3190,n0_0,q0010001_1),
       H0010001_013(h0010001_013,n3190,n0_0,q0010010_1),
       H0010010_013(h0010010_013,n3190,n0_0,q0010011_1),
       H0010011_013(h0010011_013,n3190,n0_0,q0010100_1),
       H0010100_013(h0010100_013,n3190,n0_0,q0010101_1),
       H0010101_013(h0010101_013,n3190,n0_0,q0010110_1),
       H0010110_013(h0010110_013,n3190,n0_0,q0010111_1),
       H0010111_013(h0010111_013,n3190,n0_0,q0011000_1),
       H0011000_013(h0011000_013,n3190,n0_0,q0011001_1),
       H0011001_013(h0011001_013,n3190,n0_0,q0011010_1),
       H0011010_013(h0011010_013,n3190,n0_0,q0011011_1),
       H0011011_013(h0011011_013,n3190,n0_0,q0011100_1),
       H0011100_013(h0011100_013,n3190,n0_0,q0011101_1),
       H0011101_013(h0011101_013,n3190,n0_0,q0011110_1),
       H0011110_013(h0011110_013,n3190,n0_0,q0011111_1),
       H0011111_013(h0011111_013,n3190,n0_0,q0100000_1),
       H0100000_013(h0100000_013,n3190,n0_0,q0100001_1),
       H0100001_013(h0100001_013,n3190,n0_0,q0100010_1),
       H0100010_013(h0100010_013,n3190,n0_0,q0100011_1),
       H0100011_013(h0100011_013,n3190,n0_0,q0100100_1),
       H0100100_013(h0100100_013,n3190,n0_0,q0100101_1),
       H0100101_013(h0100101_013,n3190,n0_0,q0100110_1),
       H0100110_013(h0100110_013,n3190,n0_0,q0100111_1),
       H0100111_013(h0100111_013,n3190,n0_0,q0101000_1),
       H0101000_013(h0101000_013,n3190,n0_0,q0101001_1),
       H0101001_013(h0101001_013,n3190,n0_0,q0101010_1),
       H0101010_013(h0101010_013,n3190,n0_0,q0101011_1),
       H0101011_013(h0101011_013,n3190,n0_0,q0101100_1),
       H0101100_013(h0101100_013,n3190,n0_0,q0101101_1),
       H0101101_013(h0101101_013,n3190,n0_0,q0101110_1),
       H0101110_013(h0101110_013,n3190,n0_0,q0101111_1),
       H0101111_013(h0101111_013,n3190,n0_0,q0110000_1),
       H0110000_013(h0110000_013,n3190,n0_0,q0110001_1),
       H0110001_013(h0110001_013,n3190,n0_0,q0110010_1),
       H0110010_013(h0110010_013,n3190,n0_0,q0110011_1),
       H0110011_013(h0110011_013,n3190,n0_0,q0110100_1),
       H0110100_013(h0110100_013,n3190,n0_0,q0110101_1),
       H0110101_013(h0110101_013,n3190,n0_0,q0110110_1),
       H0110110_013(h0110110_013,n3190,n0_0,q0110111_1),
       H0110111_013(h0110111_013,n3190,n0_0,q0111000_1),
       H0111000_013(h0111000_013,n3190,n0_0,q0111001_1),
       H0111001_013(h0111001_013,n3190,n0_0,q0111010_1),
       H0111010_013(h0111010_013,n3190,n0_0,q0111011_1),
       H0111011_013(h0111011_013,n3190,n0_0,q0111100_1),
       H0111100_013(h0111100_013,n3190,n0_0,q0111101_1),
       H0111101_013(h0111101_013,n3190,n0_0,q0111110_1),
       H0111110_013(h0111110_013,n3190,n0_0,q0111111_1),
       H0111111_013(h0111111_013,n3190,n0_0,q1000000_1),
       H1000000_013(h1000000_013,n3190,n0_0,q1000001_1),
       H1000001_013(h1000001_013,n3190,n0_0,q1000010_1),
       H1000010_013(h1000010_013,n3190,n0_0,q1000011_1),
       H1000011_013(h1000011_013,n3190,n0_0,q1000100_1),
       H1000100_013(h1000100_013,n3190,n0_0,q1000101_1),
       H1000101_013(h1000101_013,n3190,n0_0,q1000110_1),
       H1000110_013(h1000110_013,n3190,n0_0,q1000111_1),
       H1000111_013(h1000111_013,n3190,n0_0,q1001000_1),
       H1001000_013(h1001000_013,n3190,n0_0,q1001001_1),
       H1001001_013(h1001001_013,n3190,n0_0,q1001010_1),
       H1001010_013(h1001010_013,n3190,n0_0,q1001011_1),
       H1001011_013(h1001011_013,n3190,n0_0,q1001100_1),
       H1001100_013(h1001100_013,n3190,n0_0,q1001101_1),
       H1001101_013(h1001101_013,n3190,n0_0,q1001110_1),
       H1001110_013(h1001110_013,n3190,n0_0,q1001111_1),
       H1001111_013(h1001111_013,n3190,n0_0,q1010000_1),
       H1010000_013(h1010000_013,n3190,n0_0,q1010001_1),
       H1010001_013(h1010001_013,n3190,n0_0,q1010010_1),
       H1010010_013(h1010010_013,n3190,n0_0,q1010011_1),
       H1010011_013(h1010011_013,n3190,n0_0,q1010100_1),
       H1010100_013(h1010100_013,n3190,n0_0,q1010101_1),
       H1010101_013(h1010101_013,n3190,n0_0,q1010110_1),
       H1010110_013(h1010110_013,n3190,n0_0,q1010111_1),
       H1010111_013(h1010111_013,n3190,n0_0,q1011000_1),
       H1011000_013(h1011000_013,n3190,n0_0,q1011001_1),
       H1011001_013(h1011001_013,n3190,n0_0,q1011010_1),
       H1011010_013(h1011010_013,n3190,n0_0,q1011011_1),
       H1011011_013(h1011011_013,n3190,n0_0,q1011100_1),
       H1011100_013(h1011100_013,n3190,n0_0,q1011101_1),
       H1011101_013(h1011101_013,n3190,n0_0,q1011110_1),
       H1011110_013(h1011110_013,n3190,n0_0,q1011111_1),
       H1011111_013(h1011111_013,n3190,n0_0,q1100000_1),
       H1100000_013(h1100000_013,n3190,n0_0,q1100001_1),
       H1100001_013(h1100001_013,n3190,n0_0,q1100010_1),
       H1100010_013(h1100010_013,n3190,n0_0,q1100011_1),
       H1100011_013(h1100011_013,n3190,n0_0,q1100100_1),
       H1100100_013(h1100100_013,n3190,n0_0,q1100101_1),
       H1100101_013(h1100101_013,n3190,n0_0,q1100110_1),
       H1100110_013(h1100110_013,n3190,n0_0,q1100111_1),
       H1100111_013(h1100111_013,n3190,n0_0,q1101000_1),
       H1101000_013(h1101000_013,n3190,n0_0,q1101001_1),
       H1101001_013(h1101001_013,n3190,n0_0,q1101010_1),
       H1101010_013(h1101010_013,n3190,n0_0,q1101011_1),
       H1101011_013(h1101011_013,n3190,n0_0,q1101100_1),
       H1101100_013(h1101100_013,n3190,n0_0,q1101101_1),
       H1101101_013(h1101101_013,n3190,n0_0,q1101110_1),
       H1101110_013(h1101110_013,n3190,n0_0,q1101111_1),
       H1101111_013(h1101111_013,n3190,n0_0,q1110000_1),
       H1110000_013(h1110000_013,n3190,n0_0,q1110001_1),
       H1110001_013(h1110001_013,n3190,n0_0,q1110010_1),
       H1110010_013(h1110010_013,n3190,n0_0,q1110011_1),
       H1110011_013(h1110011_013,n3190,n0_0,q1110100_1),
       H1110100_013(h1110100_013,n3190,n0_0,q1110101_1),
       H1110101_013(h1110101_013,n3190,n0_0,q1110110_1),
       H1110110_013(h1110110_013,n3190,n0_0,q1110111_1),
       H1110111_013(h1110111_013,n3190,n0_0,q1111000_1),
       H1111000_013(h1111000_013,n3190,n0_0,q1111001_1),
       H1111001_013(h1111001_013,n3190,n0_0,q1111010_1),
       H1111010_013(h1111010_013,n3190,n0_0,q1111011_1),
       H1111011_013(h1111011_013,n3190,n0_0,q1111100_1),
       H1111100_013(h1111100_013,n3190,n0_0,q1111101_1),
       H1111101_013(h1111101_013,n3190,n0_0,q1111110_1),
       H1111110_013(h1111110_013,n3190,n0_0,q1111111_1),
       H1111111_013(h1111111_013,n3190,n0_0,dbv0);

or     H000000_0(h000000_0,h000000_011,h000000_012,h000000_013),
       H000000_1(h000000_1,h000000_111,h000000_112),
       H000001_0(h000001_0,h000001_011,h000001_012,h000001_013),
       H000001_1(h000001_1,h000001_111,h000001_112),
       H000010_0(h000010_0,h000010_011,h000010_012,h000010_013),
       H000010_1(h000010_1,h000010_111,h000010_112),
       H000011_0(h000011_0,h000011_011,h000011_012,h000011_013),
       H000011_1(h000011_1,h000011_111,h000011_112),
       H000100_0(h000100_0,h000100_011,h000100_012,h000100_013),
       H000100_1(h000100_1,h000100_111,h000100_112),
       H000101_0(h000101_0,h000101_011,h000101_012,h000101_013),
       H000101_1(h000101_1,h000101_111,h000101_112),
       H000110_0(h000110_0,h000110_011,h000110_012,h000110_013),
       H000110_1(h000110_1,h000110_111,h000110_112),
       H000111_0(h000111_0,h000111_011,h000111_012,h000111_013),
       H000111_1(h000111_1,h000111_111,h000111_112),
       H001000_0(h001000_0,h001000_011,h001000_012,h001000_013),
       H001000_1(h001000_1,h001000_111,h001000_112),
       H001001_0(h001001_0,h001001_011,h001001_012,h001001_013),
       H001001_1(h001001_1,h001001_111,h001001_112),
       H001010_0(h001010_0,h001010_011,h001010_012,h001010_013),
       H001010_1(h001010_1,h001010_111,h001010_112),
       H001011_0(h001011_0,h001011_011,h001011_012,h001011_013),
       H001011_1(h001011_1,h001011_111,h001011_112),
       H001100_0(h001100_0,h001100_011,h001100_012,h001100_013),
       H001100_1(h001100_1,h001100_111,h001100_112),
       H001101_0(h001101_0,h001101_011,h001101_012,h001101_013),
       H001101_1(h001101_1,h001101_111,h001101_112),
       H001110_0(h001110_0,h001110_011,h001110_012,h001110_013),
       H001110_1(h001110_1,h001110_111,h001110_112),
       H001111_0(h001111_0,h001111_011,h001111_012,h001111_013),
       H001111_1(h001111_1,h001111_111,h001111_112),
       H010000_0(h010000_0,h010000_011,h010000_012,h010000_013),
       H010000_1(h010000_1,h010000_111,h010000_112),
       H010001_0(h010001_0,h010001_011,h010001_012,h010001_013),
       H010001_1(h010001_1,h010001_111,h010001_112),
       H010010_0(h010010_0,h010010_011,h010010_012,h010010_013),
       H010010_1(h010010_1,h010010_111,h010010_112),
       H010011_0(h010011_0,h010011_011,h010011_012,h010011_013),
       H010011_1(h010011_1,h010011_111,h010011_112),
       H010100_0(h010100_0,h010100_011,h010100_012,h010100_013),
       H010100_1(h010100_1,h010100_111,h010100_112),
       H010101_0(h010101_0,h010101_011,h010101_012,h010101_013),
       H010101_1(h010101_1,h010101_111,h010101_112),
       H010110_0(h010110_0,h010110_011,h010110_012,h010110_013),
       H010110_1(h010110_1,h010110_111,h010110_112),
       H010111_0(h010111_0,h010111_011,h010111_012,h010111_013),
       H010111_1(h010111_1,h010111_111,h010111_112),
       H011000_0(h011000_0,h011000_011,h011000_012,h011000_013),
       H011000_1(h011000_1,h011000_111,h011000_112),
       H011001_0(h011001_0,h011001_011,h011001_012,h011001_013),
       H011001_1(h011001_1,h011001_111,h011001_112),
       H011010_0(h011010_0,h011010_011,h011010_012,h011010_013),
       H011010_1(h011010_1,h011010_111,h011010_112),
       H011011_0(h011011_0,h011011_011,h011011_012,h011011_013),
       H011011_1(h011011_1,h011011_111,h011011_112),
       H011100_0(h011100_0,h011100_011,h011100_012,h011100_013),
       H011100_1(h011100_1,h011100_111,h011100_112),
       H011101_0(h011101_0,h011101_011,h011101_012,h011101_013),
       H011101_1(h011101_1,h011101_111,h011101_112),
       H011110_0(h011110_0,h011110_011,h011110_012,h011110_013,q11_1),
       H011110_1(h011110_1,h011110_111,h011110_112,q11_1),
       H011111_0(h011111_0,h011111_011,h011111_012,h011111_013,q11_1),
       H011111_1(h011111_1,h011111_111,h011111_112,q11_1),
       H100000_0(h100000_0,h100000_011,h100000_012,h100000_013,q11_1),
       H100000_1(h100000_1,h100000_111,h100000_112,q11_1),
       H100001_0(h100001_0,h100001_011,h100001_012,h100001_013,q11_1),
       H100001_1(h100001_1,h100001_111,h100001_112,q11_1),
       H100010_0(h100010_0,h100010_011,h100010_012,h100010_013),
       H100010_1(h100010_1,h100010_111,h100010_112),
       H100011_0(h100011_0,h100011_011,h100011_012,h100011_013),
       H100011_1(h100011_1,h100011_111,h100011_112),
       H100100_0(h100100_0,h100100_011,h100100_012,h100100_013),
       H100100_1(h100100_1,h100100_111,h100100_112),
       H100101_0(h100101_0,h100101_011,h100101_012,h100101_013),
       H100101_1(h100101_1,h100101_111,h100101_112),
       H100110_0(h100110_0,h100110_011,h100110_012,h100110_013),
       H100110_1(h100110_1,h100110_111,h100110_112),
       H100111_0(h100111_0,h100111_011,h100111_012,h100111_013),
       H100111_1(h100111_1,h100111_111,h100111_112),
       H101000_0(h101000_0,h101000_011,h101000_012,h101000_013),
       H101000_1(h101000_1,h101000_111,h101000_112),
       H101001_0(h101001_0,h101001_011,h101001_012,h101001_013),
       H101001_1(h101001_1,h101001_111,h101001_112),
       H101010_0(h101010_0,h101010_011,h101010_012,h101010_013),
       H101010_1(h101010_1,h101010_111,h101010_112),
       H101011_0(h101011_0,h101011_011,h101011_012,h101011_013),
       H101011_1(h101011_1,h101011_111,h101011_112),
       H101100_0(h101100_0,h101100_011,h101100_012,h101100_013),
       H101100_1(h101100_1,h101100_111,h101100_112),
       H101101_0(h101101_0,h101101_011,h101101_012,h101101_013),
       H101101_1(h101101_1,h101101_111,h101101_112),
       H101110_0(h101110_0,h101110_011,h101110_012,h101110_013),
       H101110_1(h101110_1,h101110_111,h101110_112),
       H101111_0(h101111_0,h101111_011,h101111_012,h101111_013),
       H101111_1(h101111_1,h101111_111,h101111_112),
       H110000_0(h110000_0,h110000_011,h110000_012,h110000_013),
       H110000_1(h110000_1,h110000_111,h110000_112),
       H110001_0(h110001_0,h110001_011,h110001_012,h110001_013),
       H110001_1(h110001_1,h110001_111,h110001_112),
       H110010_0(h110010_0,h110010_011,h110010_012,h110010_013),
       H110010_1(h110010_1,h110010_111,h110010_112),
       H110011_0(h110011_0,h110011_011,h110011_012,h110011_013),
       H110011_1(h110011_1,h110011_111,h110011_112),
       H110100_0(h110100_0,h110100_011,h110100_012,h110100_013),
       H110100_1(h110100_1,h110100_111,h110100_112),
       H110101_0(h110101_0,h110101_011,h110101_012,h110101_013),
       H110101_1(h110101_1,h110101_111,h110101_112),
       H110110_0(h110110_0,h110110_011,h110110_012,h110110_013),
       H110110_1(h110110_1,h110110_111,h110110_112),
       H110111_0(h110111_0,h110111_011,h110111_012,h110111_013),
       H110111_1(h110111_1,h110111_111,h110111_112),
       H111000_0(h111000_0,h111000_011,h111000_012,h111000_013),
       H111000_1(h111000_1,h111000_111,h111000_112),
       H111001_0(h111001_0,h111001_011,h111001_012,h111001_013),
       H111001_1(h111001_1,h111001_111,h111001_112),
       H111010_0(h111010_0,h111010_011,h111010_012,h111010_013),
       H111010_1(h111010_1,h111010_111,h111010_112),
       H111011_0(h111011_0,h111011_011,h111011_012,h111011_013),
       H111011_1(h111011_1,h111011_111,h111011_112),
       H111100_0(h111100_0,h111100_011,h111100_012,h111100_013),
       H111100_1(h111100_1,h111100_111,h111100_112),
       H111101_0(h111101_0,h111101_011,h111101_012,h111101_013),
       H111101_1(h111101_1,h111101_111,h111101_112),
       H111110_0(h111110_0,h111110_011,h111110_012,h111110_013),
       H111110_1(h111110_1,h111110_111,h111110_112),
       H111111_0(h111111_0,h111111_011,h111111_012,h111111_013),
       H111111_1(h111111_1,h111111_111,h111111_112);

and    H000000_011(h000000_011,o9150,q000000_0),
       H000000_111(h000000_111,o9150,q000000_0),
       H000001_011(h000001_011,o9150,q000001_0),
       H000001_111(h000001_111,o9150,q000001_0),
       H000010_011(h000010_011,o9150,q000010_0,n11_1),
       H000010_111(h000010_111,o9150,q000010_0,n11_1),
       H000011_011(h000011_011,o9150,q000011_0,n11_1),
       H000011_111(h000011_111,o9150,q000011_0,n11_1),
       H000100_011(h000100_011,o9150,q000100_0,n11_1),
       H000100_111(h000100_111,o9150,q000100_0,n11_1),
       H000101_011(h000101_011,o9150,q000101_0,n11_1),
       H000101_111(h000101_111,o9150,q000101_0,n11_1),
       H000110_011(h000110_011,o9150,q000110_0,n11_1),
       H000110_111(h000110_111,o9150,q000110_0,n11_1),
       H000111_011(h000111_011,o9150,q000111_0,n11_1),
       H000111_111(h000111_111,o9150,q000111_0,n11_1),
       H001000_011(h001000_011,o9150,q001000_0,n11_1),
       H001000_111(h001000_111,o9150,q001000_0,n11_1),
       H001001_011(h001001_011,o9150,q001001_0,n11_1),
       H001001_111(h001001_111,o9150,q001001_0,n11_1),
       H001010_011(h001010_011,o9150,q001010_0,n11_1),
       H001010_111(h001010_111,o9150,q001010_0,n11_1),
       H001011_011(h001011_011,o9150,q001011_0,n11_1),
       H001011_111(h001011_111,o9150,q001011_0,n11_1),
       H001100_011(h001100_011,o9150,q001100_0,n11_1),
       H001100_111(h001100_111,o9150,q001100_0,n11_1),
       H001101_011(h001101_011,o9150,q001101_0,n11_1),
       H001101_111(h001101_111,o9150,q001101_0,n11_1),
       H001110_011(h001110_011,o9150,q001110_0,n11_1),
       H001110_111(h001110_111,o9150,q001110_0,n11_1),
       H001111_011(h001111_011,o9150,q001111_0,n11_1),
       H001111_111(h001111_111,o9150,q001111_0,n11_1),
       H010000_011(h010000_011,o9150,q010000_0,n11_1),
       H010000_111(h010000_111,o9150,q010000_0,n11_1),
       H010001_011(h010001_011,o9150,q010001_0,n11_1),
       H010001_111(h010001_111,o9150,q010001_0,n11_1),
       H010010_011(h010010_011,o9150,q010010_0,n11_1),
       H010010_111(h010010_111,o9150,q010010_0,n11_1),
       H010011_011(h010011_011,o9150,q010011_0,n11_1),
       H010011_111(h010011_111,o9150,q010011_0,n11_1),
       H010100_011(h010100_011,o9150,q010100_0,n11_1),
       H010100_111(h010100_111,o9150,q010100_0,n11_1),
       H010101_011(h010101_011,o9150,q010101_0,n11_1),
       H010101_111(h010101_111,o9150,q010101_0,n11_1),
       H010110_011(h010110_011,o9150,q010110_0,n11_1),
       H010110_111(h010110_111,o9150,q010110_0,n11_1),
       H010111_011(h010111_011,o9150,q010111_0,n11_1),
       H010111_111(h010111_111,o9150,q010111_0,n11_1),
       H011000_011(h011000_011,o9150,q011000_0,n11_1),
       H011000_111(h011000_111,o9150,q011000_0,n11_1),
       H011001_011(h011001_011,o9150,q011001_0,n11_1),
       H011001_111(h011001_111,o9150,q011001_0,n11_1),
       H011010_011(h011010_011,o9150,q011010_0,n11_1),
       H011010_111(h011010_111,o9150,q011010_0,n11_1),
       H011011_011(h011011_011,o9150,q011011_0,n11_1),
       H011011_111(h011011_111,o9150,q011011_0,n11_1),
       H011100_011(h011100_011,o9150,q011100_0,n11_1),
       H011100_111(h011100_111,o9150,q011100_0,n11_1),
       H011101_011(h011101_011,o9150,q011101_0,n11_1),
       H011101_111(h011101_111,o9150,q011101_0,n11_1),
       H011110_011(h011110_011,o9150,q011110_0,n11_1),
       H011110_111(h011110_111,o9150,q011110_0,n11_1),
       H011111_011(h011111_011,o9150,q011111_0,n11_1),
       H011111_111(h011111_111,o9150,q011111_0,n11_1),
       H100000_011(h100000_011,o9150,q100000_0,n11_1),
       H100000_111(h100000_111,o9150,q100000_0,n11_1),
       H100001_011(h100001_011,o9150,q100001_0,n11_1),
       H100001_111(h100001_111,o9150,q100001_0,n11_1),
       H100010_011(h100010_011,o9150,q100010_0,n11_1),
       H100010_111(h100010_111,o9150,q100010_0,n11_1),
       H100011_011(h100011_011,o9150,q100011_0,n11_1),
       H100011_111(h100011_111,o9150,q100011_0,n11_1),
       H100100_011(h100100_011,o9150,q100100_0,n11_1),
       H100100_111(h100100_111,o9150,q100100_0,n11_1),
       H100101_011(h100101_011,o9150,q100101_0,n11_1),
       H100101_111(h100101_111,o9150,q100101_0,n11_1),
       H100110_011(h100110_011,o9150,q100110_0,n11_1),
       H100110_111(h100110_111,o9150,q100110_0,n11_1),
       H100111_011(h100111_011,o9150,q100111_0,n11_1),
       H100111_111(h100111_111,o9150,q100111_0,n11_1),
       H101000_011(h101000_011,o9150,q101000_0,n11_1),
       H101000_111(h101000_111,o9150,q101000_0,n11_1),
       H101001_011(h101001_011,o9150,q101001_0,n11_1),
       H101001_111(h101001_111,o9150,q101001_0,n11_1),
       H101010_011(h101010_011,o9150,q101010_0,n11_1),
       H101010_111(h101010_111,o9150,q101010_0,n11_1),
       H101011_011(h101011_011,o9150,q101011_0,n11_1),
       H101011_111(h101011_111,o9150,q101011_0,n11_1),
       H101100_011(h101100_011,o9150,q101100_0,n11_1),
       H101100_111(h101100_111,o9150,q101100_0,n11_1),
       H101101_011(h101101_011,o9150,q101101_0,n11_1),
       H101101_111(h101101_111,o9150,q101101_0,n11_1),
       H101110_011(h101110_011,o9150,q101110_0,n11_1),
       H101110_111(h101110_111,o9150,q101110_0,n11_1),
       H101111_011(h101111_011,o9150,q101111_0,n11_1),
       H101111_111(h101111_111,o9150,q101111_0,n11_1),
       H110000_011(h110000_011,o9150,q110000_0,n11_1),
       H110000_111(h110000_111,o9150,q110000_0,n11_1),
       H110001_011(h110001_011,o9150,q110001_0,n11_1),
       H110001_111(h110001_111,o9150,q110001_0,n11_1),
       H110010_011(h110010_011,o9150,q110010_0,n11_1),
       H110010_111(h110010_111,o9150,q110010_0,n11_1),
       H110011_011(h110011_011,o9150,q110011_0,n11_1),
       H110011_111(h110011_111,o9150,q110011_0,n11_1),
       H110100_011(h110100_011,o9150,q110100_0,n11_1),
       H110100_111(h110100_111,o9150,q110100_0,n11_1),
       H110101_011(h110101_011,o9150,q110101_0,n11_1),
       H110101_111(h110101_111,o9150,q110101_0,n11_1),
       H110110_011(h110110_011,o9150,q110110_0,n11_1),
       H110110_111(h110110_111,o9150,q110110_0,n11_1),
       H110111_011(h110111_011,o9150,q110111_0,n11_1),
       H110111_111(h110111_111,o9150,q110111_0,n11_1),
       H111000_011(h111000_011,o9150,q111000_0,n11_1),
       H111000_111(h111000_111,o9150,q111000_0,n11_1),
       H111001_011(h111001_011,o9150,q111001_0,n11_1),
       H111001_111(h111001_111,o9150,q111001_0,n11_1),
       H111010_011(h111010_011,o9150,q111010_0,n11_1),
       H111010_111(h111010_111,o9150,q111010_0,n11_1),
       H111011_011(h111011_011,o9150,q111011_0,n11_1),
       H111011_111(h111011_111,o9150,q111011_0,n11_1),
       H111100_011(h111100_011,o9150,q111100_0,n11_1),
       H111100_111(h111100_111,o9150,q111100_0,n11_1),
       H111101_011(h111101_011,o9150,q111101_0,n11_1),
       H111101_111(h111101_111,o9150,q111101_0,n11_1),
       H111110_011(h111110_011,o9150,q111110_0),
       H111110_111(h111110_111,o9150,q111110_0),
       H111111_011(h111111_011,o9150,q111111_0),
       H111111_111(h111111_111,o9150,q111111_0),
       H000000_012(h000000_012,n9150,q1_0,q000000_1),
       H000000_112(h000000_112,n9150,q000000_1),
       H000001_012(h000001_012,n9150,q1_0,q000001_1),
       H000001_112(h000001_112,n9150,q000001_1),
       H000010_012(h000010_012,n9150,q1_0,dbv0),
       H000010_112(h000010_112,n9150,q000010_1),
       H000011_012(h000011_012,n9150,q1_0,q000010_1),
       H000011_112(h000011_112,n9150,q000011_1),
       H000100_012(h000100_012,n9150,q1_0,q000011_1),
       H000100_112(h000100_112,n9150,q000100_1),
       H000101_012(h000101_012,n9150,q1_0,q000100_1),
       H000101_112(h000101_112,n9150,q000101_1),
       H000110_012(h000110_012,n9150,q1_0,q000101_1),
       H000110_112(h000110_112,n9150,q000110_1),
       H000111_012(h000111_012,n9150,q1_0,q000110_1),
       H000111_112(h000111_112,n9150,q000111_1),
       H001000_012(h001000_012,n9150,q1_0,q000111_1),
       H001000_112(h001000_112,n9150,q001000_1),
       H001001_012(h001001_012,n9150,q1_0,q001000_1),
       H001001_112(h001001_112,n9150,q001001_1),
       H001010_012(h001010_012,n9150,q1_0,q001001_1),
       H001010_112(h001010_112,n9150,q001010_1),
       H001011_012(h001011_012,n9150,q1_0,q001010_1),
       H001011_112(h001011_112,n9150,q001011_1),
       H001100_012(h001100_012,n9150,q1_0,q001011_1),
       H001100_112(h001100_112,n9150,q001100_1),
       H001101_012(h001101_012,n9150,q1_0,q001100_1),
       H001101_112(h001101_112,n9150,q001101_1),
       H001110_012(h001110_012,n9150,q1_0,q001101_1),
       H001110_112(h001110_112,n9150,q001110_1),
       H001111_012(h001111_012,n9150,q1_0,q001110_1),
       H001111_112(h001111_112,n9150,q001111_1),
       H010000_012(h010000_012,n9150,q1_0,q001111_1),
       H010000_112(h010000_112,n9150,q010000_1),
       H010001_012(h010001_012,n9150,q1_0,q010000_1),
       H010001_112(h010001_112,n9150,q010001_1),
       H010010_012(h010010_012,n9150,q1_0,q010001_1),
       H010010_112(h010010_112,n9150,q010010_1),
       H010011_012(h010011_012,n9150,q1_0,q010010_1),
       H010011_112(h010011_112,n9150,q010011_1),
       H010100_012(h010100_012,n9150,q1_0,q010011_1),
       H010100_112(h010100_112,n9150,q010100_1),
       H010101_012(h010101_012,n9150,q1_0,q010100_1),
       H010101_112(h010101_112,n9150,q010101_1),
       H010110_012(h010110_012,n9150,q1_0,q010101_1),
       H010110_112(h010110_112,n9150,q010110_1),
       H010111_012(h010111_012,n9150,q1_0,q010110_1),
       H010111_112(h010111_112,n9150,q010111_1),
       H011000_012(h011000_012,n9150,q1_0,q010111_1),
       H011000_112(h011000_112,n9150,q011000_1),
       H011001_012(h011001_012,n9150,q1_0,q011000_1),
       H011001_112(h011001_112,n9150,q011001_1),
       H011010_012(h011010_012,n9150,q1_0,q011001_1),
       H011010_112(h011010_112,n9150,q011010_1),
       H011011_012(h011011_012,n9150,q1_0,q011010_1),
       H011011_112(h011011_112,n9150,q011011_1),
       H011100_012(h011100_012,n9150,q1_0,q011011_1),
       H011100_112(h011100_112,n9150,q011100_1),
       H011101_012(h011101_012,n9150,q1_0,q011100_1),
       H011101_112(h011101_112,n9150,q011101_1),
       H011110_012(h011110_012,n9150,q1_0,q011101_1),
       H011110_112(h011110_112,n9150,q011110_1),
       H011111_012(h011111_012,n9150,q1_0,q011110_1),
       H011111_112(h011111_112,n9150,q011111_1),
       H100000_012(h100000_012,n9150,q1_0,q011111_1),
       H100000_112(h100000_112,n9150,q100000_1),
       H100001_012(h100001_012,n9150,q1_0,q100000_1),
       H100001_112(h100001_112,n9150,q100001_1),
       H100010_012(h100010_012,n9150,q1_0,q100001_1),
       H100010_112(h100010_112,n9150,q100010_1),
       H100011_012(h100011_012,n9150,q1_0,q100010_1),
       H100011_112(h100011_112,n9150,q100011_1),
       H100100_012(h100100_012,n9150,q1_0,q100011_1),
       H100100_112(h100100_112,n9150,q100100_1),
       H100101_012(h100101_012,n9150,q1_0,q100100_1),
       H100101_112(h100101_112,n9150,q100101_1),
       H100110_012(h100110_012,n9150,q1_0,q100101_1),
       H100110_112(h100110_112,n9150,q100110_1),
       H100111_012(h100111_012,n9150,q1_0,q100110_1),
       H100111_112(h100111_112,n9150,q100111_1),
       H101000_012(h101000_012,n9150,q1_0,q100111_1),
       H101000_112(h101000_112,n9150,q101000_1),
       H101001_012(h101001_012,n9150,q1_0,q101000_1),
       H101001_112(h101001_112,n9150,q101001_1),
       H101010_012(h101010_012,n9150,q1_0,q101001_1),
       H101010_112(h101010_112,n9150,q101010_1),
       H101011_012(h101011_012,n9150,q1_0,q101010_1),
       H101011_112(h101011_112,n9150,q101011_1),
       H101100_012(h101100_012,n9150,q1_0,q101011_1),
       H101100_112(h101100_112,n9150,q101100_1),
       H101101_012(h101101_012,n9150,q1_0,q101100_1),
       H101101_112(h101101_112,n9150,q101101_1),
       H101110_012(h101110_012,n9150,q1_0,q101101_1),
       H101110_112(h101110_112,n9150,q101110_1),
       H101111_012(h101111_012,n9150,q1_0,q101110_1),
       H101111_112(h101111_112,n9150,q101111_1),
       H110000_012(h110000_012,n9150,q1_0,q101111_1),
       H110000_112(h110000_112,n9150,q110000_1),
       H110001_012(h110001_012,n9150,q1_0,q110000_1),
       H110001_112(h110001_112,n9150,q110001_1),
       H110010_012(h110010_012,n9150,q1_0,q110001_1),
       H110010_112(h110010_112,n9150,q110010_1),
       H110011_012(h110011_012,n9150,q1_0,q110010_1),
       H110011_112(h110011_112,n9150,q110011_1),
       H110100_012(h110100_012,n9150,q1_0,q110011_1),
       H110100_112(h110100_112,n9150,q110100_1),
       H110101_012(h110101_012,n9150,q1_0,q110100_1),
       H110101_112(h110101_112,n9150,q110101_1),
       H110110_012(h110110_012,n9150,q1_0,q110101_1),
       H110110_112(h110110_112,n9150,q110110_1),
       H110111_012(h110111_012,n9150,q1_0,q110110_1),
       H110111_112(h110111_112,n9150,q110111_1),
       H111000_012(h111000_012,n9150,q1_0,q110111_1),
       H111000_112(h111000_112,n9150,q111000_1),
       H111001_012(h111001_012,n9150,q1_0,q111000_1),
       H111001_112(h111001_112,n9150,q111001_1),
       H111010_012(h111010_012,n9150,q1_0,q111001_1),
       H111010_112(h111010_112,n9150,q111010_1),
       H111011_012(h111011_012,n9150,q1_0,q111010_1),
       H111011_112(h111011_112,n9150,q111011_1),
       H111100_012(h111100_012,n9150,q1_0,q111011_1),
       H111100_112(h111100_112,n9150,q111100_1),
       H111101_012(h111101_012,n9150,q1_0,q111100_1),
       H111101_112(h111101_112,n9150,q111101_1),
       H111110_012(h111110_012,n9150,q1_0,q111110_1),
       H111110_112(h111110_112,n9150,q111110_1),
       H111111_012(h111111_012,n9150,q1_0,q111111_1),
       H111111_112(h111111_112,n9150,q111111_1),
       H000000_013(h000000_013,n9150,n1_0,q000000_1),
       H000001_013(h000001_013,n9150,n1_0,q000001_1),
       H000010_013(h000010_013,n9150,n1_0,q000011_1),
       H000011_013(h000011_013,n9150,n1_0,q000100_1),
       H000100_013(h000100_013,n9150,n1_0,q000101_1),
       H000101_013(h000101_013,n9150,n1_0,q000110_1),
       H000110_013(h000110_013,n9150,n1_0,q000111_1),
       H000111_013(h000111_013,n9150,n1_0,q001000_1),
       H001000_013(h001000_013,n9150,n1_0,q001001_1),
       H001001_013(h001001_013,n9150,n1_0,q001010_1),
       H001010_013(h001010_013,n9150,n1_0,q001011_1),
       H001011_013(h001011_013,n9150,n1_0,q001100_1),
       H001100_013(h001100_013,n9150,n1_0,q001101_1),
       H001101_013(h001101_013,n9150,n1_0,q001110_1),
       H001110_013(h001110_013,n9150,n1_0,q001111_1),
       H001111_013(h001111_013,n9150,n1_0,q010000_1),
       H010000_013(h010000_013,n9150,n1_0,q010001_1),
       H010001_013(h010001_013,n9150,n1_0,q010010_1),
       H010010_013(h010010_013,n9150,n1_0,q010011_1),
       H010011_013(h010011_013,n9150,n1_0,q010100_1),
       H010100_013(h010100_013,n9150,n1_0,q010101_1),
       H010101_013(h010101_013,n9150,n1_0,q010110_1),
       H010110_013(h010110_013,n9150,n1_0,q010111_1),
       H010111_013(h010111_013,n9150,n1_0,q011000_1),
       H011000_013(h011000_013,n9150,n1_0,q011001_1),
       H011001_013(h011001_013,n9150,n1_0,q011010_1),
       H011010_013(h011010_013,n9150,n1_0,q011011_1),
       H011011_013(h011011_013,n9150,n1_0,q011100_1),
       H011100_013(h011100_013,n9150,n1_0,q011101_1),
       H011101_013(h011101_013,n9150,n1_0,q011110_1),
       H011110_013(h011110_013,n9150,n1_0,q011111_1),
       H011111_013(h011111_013,n9150,n1_0,q100000_1),
       H100000_013(h100000_013,n9150,n1_0,q100001_1),
       H100001_013(h100001_013,n9150,n1_0,q100010_1),
       H100010_013(h100010_013,n9150,n1_0,q100011_1),
       H100011_013(h100011_013,n9150,n1_0,q100100_1),
       H100100_013(h100100_013,n9150,n1_0,q100101_1),
       H100101_013(h100101_013,n9150,n1_0,q100110_1),
       H100110_013(h100110_013,n9150,n1_0,q100111_1),
       H100111_013(h100111_013,n9150,n1_0,q101000_1),
       H101000_013(h101000_013,n9150,n1_0,q101001_1),
       H101001_013(h101001_013,n9150,n1_0,q101010_1),
       H101010_013(h101010_013,n9150,n1_0,q101011_1),
       H101011_013(h101011_013,n9150,n1_0,q101100_1),
       H101100_013(h101100_013,n9150,n1_0,q101101_1),
       H101101_013(h101101_013,n9150,n1_0,q101110_1),
       H101110_013(h101110_013,n9150,n1_0,q101111_1),
       H101111_013(h101111_013,n9150,n1_0,q110000_1),
       H110000_013(h110000_013,n9150,n1_0,q110001_1),
       H110001_013(h110001_013,n9150,n1_0,q110010_1),
       H110010_013(h110010_013,n9150,n1_0,q110011_1),
       H110011_013(h110011_013,n9150,n1_0,q110100_1),
       H110100_013(h110100_013,n9150,n1_0,q110101_1),
       H110101_013(h110101_013,n9150,n1_0,q110110_1),
       H110110_013(h110110_013,n9150,n1_0,q110111_1),
       H110111_013(h110111_013,n9150,n1_0,q111000_1),
       H111000_013(h111000_013,n9150,n1_0,q111001_1),
       H111001_013(h111001_013,n9150,n1_0,q111010_1),
       H111010_013(h111010_013,n9150,n1_0,q111011_1),
       H111011_013(h111011_013,n9150,n1_0,q111100_1),
       H111100_013(h111100_013,n9150,n1_0,q111101_1),
       H111101_013(h111101_013,n9150,n1_0,dbv0),
       H111110_013(h111110_013,n9150,n1_0,q111110_1),
       H111111_013(h111111_013,n9150,n1_0,q111111_1);

not    N0001(n0001,q0001);
xor    X0002(x0002,q0002,q0001),
       X0003(x0003,q0003,a0003),
       X0004(x0004,q0004,a0004),
       X0005(x0005,q0005,a0005),
       X0006(x0006,q0006,a0006),
       X0007(x0007,q0007,a0007),
       X0008(x0008,q0008,a0008),
       X0009(x0009,q0009,a0009),
       X0010(x0010,q0010,a0010),
       X0011(x0011,q0011,a0011),
       X0012(x0012,q0012,a0012),
       X0013(x0013,q0013,a0013),
       X0014(x0014,q0014,a0014),
       X0015(x0015,q0015,a0015),
       X0016(x0016,q0016,a0016),
       X0017(x0017,q0017,a0017),
       X0018(x0018,q0018,a0018),
       X0019(x0019,q0019,a0019),
       X0020(x0020,q0020,a0020),
       X0021(x0021,q0021,a0021),
       X0022(x0022,q0022,a0022),
       X0023(x0023,q0023,a0023),
       X0024(x0024,q0024,a0024),
       X0025(x0025,q0025,a0025),
       X0026(x0026,q0026,a0026),
       X0027(x0027,q0027,a0027),
       X0028(x0028,q0028,a0028),
       X0029(x0029,q0029,a0029),
       X0030(x0030,q0030,a0030);

and    A0003(a0003,q0002,q0001),
       A0004(a0004,a0003,q0003),
       A0005(a0005,a0004,q0004),
       A0006(a0006,a0005,q0005),
       A0007(a0007,a0006,q0006),
       A0008(a0008,a0007,q0007),
       A0009(a0009,a0008,q0008),
       A0010(a0010,a0009,q0009),
       A0011(a0011,a0010,q0010),
       A0012(a0012,a0011,q0011),
       A0013(a0013,a0012,q0012),
       A0014(a0014,a0013,q0013),
       A0015(a0015,a0014,q0014),
       A0016(a0016,a0015,q0015),
       A0017(a0017,a0016,q0016),
       A0018(a0018,a0017,q0017),
       A0019(a0019,a0018,q0018),
       A0020(a0020,a0019,q0019),
       A0021(a0021,a0020,q0020),
       A0022(a0022,a0021,q0021),
       A0023(a0023,a0022,q0022),
       A0024(a0024,a0023,q0023),
       A0025(a0025,a0024,q0024),
       A0026(a0026,a0025,q0025),
       A0027(a0027,a0026,q0026),
       A0028(a0028,a0027,q0027),
       A0029(a0029,a0028,q0028),
       A0030(a0030,a0029,q0029);
//x
not    N0031(n0031,q0031);
xor    X0032(x0032,q0032,q0031),
       X0033(x0033,q0033,a0033),
       X0034(x0034,q0034,a0034),
       X0035(x0035,q0035,a0035),
       X0036(x0036,q0036,a0036),
       X0037(x0037,q0037,a0037),
       X0038(x0038,q0038,a0038),
       X0039(x0039,q0039,a0039),
       X0040(x0040,q0040,a0040),
       X0041(x0041,q0041,a0041),
       X0042(x0042,q0042,a0042),
       X0043(x0043,q0043,a0043),
       X0044(x0044,q0044,a0044),
       X0045(x0045,q0045,a0045),
       X0046(x0046,q0046,a0046),
       X0047(x0047,q0047,a0047),
       X0048(x0048,q0048,a0048),
       X0049(x0049,q0049,a0049),
       X0050(x0050,q0050,a0050),
       X0051(x0051,q0051,a0051),
       X0052(x0052,q0052,a0052),
       X0053(x0053,q0053,a0053),
       X0054(x0054,q0054,a0054),
       X0055(x0055,q0055,a0055),
       X0056(x0056,q0056,a0056),
       X0057(x0057,q0057,a0057),
       X0058(x0058,q0058,a0058),
       X0059(x0059,q0059,a0059),
       X0060(x0060,q0060,a0060);

and    A0033(a0033,q0032,q0031),
       A0034(a0034,a0033,q0033),
       A0035(a0035,a0034,q0034),
       A0036(a0036,a0035,q0035),
       A0037(a0037,a0036,q0036),
       A0038(a0038,a0037,q0037),
       A0039(a0039,a0038,q0038),
       A0040(a0040,a0039,q0039),
       A0041(a0041,a0040,q0040),
       A0042(a0042,a0041,q0041),
       A0043(a0043,a0042,q0042),
       A0044(a0044,a0043,q0043),
       A0045(a0045,a0044,q0044),
       A0046(a0046,a0045,q0045),
       A0047(a0047,a0046,q0046),
       A0048(a0048,a0047,q0047),
       A0049(a0049,a0048,q0048),
       A0050(a0050,a0049,q0049),
       A0051(a0051,a0050,q0050),
       A0052(a0052,a0051,q0051),
       A0053(a0053,a0052,q0052),
       A0054(a0054,a0053,q0053),
       A0055(a0055,a0054,q0054),
       A0056(a0056,a0055,q0055),
       A0057(a0057,a0056,q0056),
       A0058(a0058,a0057,q0057),
       A0059(a0059,a0058,q0058),
       A0060(a0060,a0059,q0059);

xor    X0061(x0061,q0061,q0031),
       X0062(x0062,q0062,q0032),
       X0063(x0063,q0063,q0033),
       X0064(x0064,q0064,q0034),
       X0065(x0065,q0065,q0035),
       X0066(x0066,q0066,q0036),
       X0067(x0067,q0067,q0037),
       X0068(x0068,q0068,q0038),
       X0069(x0069,q0069,q0039),
       X0070(x0070,q0070,q0040),
       X0071(x0071,q0071,q0041),
       X0072(x0072,q0072,q0042),
       X0073(x0073,q0073,q0043),
       X0074(x0074,q0074,q0044),
       X0075(x0075,q0075,q0045),
       X0076(x0076,q0076,q0046),
       X0077(x0077,q0077,q0047),
       X0078(x0078,q0078,q0048),
       X0079(x0079,q0079,q0049),
       X0080(x0080,q0080,q0050),
       X0081(x0081,q0081,q0051),
       X0082(x0082,q0082,q0052),
       X0083(x0083,q0083,q0053),
       X0084(x0084,q0084,q0054),
       X0085(x0085,q0085,q0055),
       X0086(x0086,q0086,q0056),
       X0087(x0087,q0087,q0057),
       X0088(x0088,q0088,q0058),
       X0089(x0089,q0089,q0059),
       X0090(x0090,q0090,q0060);

and    A0061(a0061,n0031,o3190,n11_1),
       A0062(a0062,x0032,o3190,n11_1),
       A0063(a0063,x0033,o3190,n11_1),
       A0064(a0064,x0034,o3190,n11_1),
       A0065(a0065,x0035,o3190,n11_1),
       A0066(a0066,x0036,o3190,n11_1),
       A0067(a0067,x0037,o3190,n11_1),
       A0068(a0068,x0038,o3190,n11_1),
       A0069(a0069,x0039,o3190,n11_1),
       A0070(a0070,x0040,o3190,n11_1),
       A0071(a0071,x0041,o3190,n11_1),
       A0072(a0072,x0042,o3190,n11_1),
       A0073(a0073,x0043,o3190,n11_1),
       A0074(a0074,x0044,o3190,n11_1),
       A0075(a0075,x0045,o3190,n11_1),
       A0076(a0076,x0046,o3190,n11_1),
       A0077(a0077,x0047,o3190,n11_1),
       A0078(a0078,x0048,o3190,n11_1),
       A0079(a0079,x0049,o3190,n11_1),
       A0080(a0080,x0050,o3190,n11_1),
       A0081(a0081,x0051,o3190,n11_1),
       A0082(a0082,x0052,o3190,n11_1),
       A0083(a0083,x0053,o3190,n11_1),
       A0084(a0084,x0054,o3190,n11_1),
       A0085(a0085,x0055,o3190,n11_1),
       A0086(a0086,x0056,o3190,n11_1),
       A0087(a0087,x0057,o3190,n11_1),
       A0088(a0088,x0058,o3190,n11_1),
       A0089(a0089,x0059,o3190,n11_1),
       A0090(a0090,x0060,o3190,n11_1);

or     H006101(h006101,h006111,h006112),
       H006102(h006102,dbv0,dbv0),
       H006201(h006201,h006211,h006212),
       H006202(h006202,dbv0,dbv0),
       H006301(h006301,h006311,h006312),
       H006302(h006302,dbv0,dbv0),
       H006401(h006401,h006411,h006412),
       H006402(h006402,dbv0,dbv0),
       H006501(h006501,h006511,h006512),
       H006502(h006502,dbv0,dbv0),
       H006601(h006601,h006611,h006612),
       H006602(h006602,dbv0,dbv0),
       H006701(h006701,h006711,h006712),
       H006702(h006702,dbv0,dbv0),
       H006801(h006801,h006811,h006812),
       H006802(h006802,dbv0,dbv0),
       H006901(h006901,h006911,h006912),
       H006902(h006902,dbv0,dbv0),
       H007001(h007001,h007011,h007012),
       H007002(h007002,dbv0,dbv0),
       H007101(h007101,h007111,h007112),
       H007102(h007102,dbv0,dbv0),
       H007201(h007201,h007211,h007212),
       H007202(h007202,dbv0,dbv0),
       H007301(h007301,h007311,h007312),
       H007302(h007302,dbv0,dbv0),
       H007401(h007401,h007411,h007412),
       H007402(h007402,dbv0,dbv0),
       H007501(h007501,h007511,h007512),
       H007502(h007502,dbv0,dbv0),
       H007601(h007601,h007611,h007612),
       H007602(h007602,dbv0,dbv0),
       H007701(h007701,h007711,h007712),
       H007702(h007702,dbv0,dbv0),
       H007801(h007801,h007811,h007812),
       H007802(h007802,dbv0,dbv0),
       H007901(h007901,h007911,h007912),
       H007902(h007902,dbv0,dbv0),
       H008001(h008001,h008011,h008012),
       H008002(h008002,dbv0,dbv0),
       H008101(h008101,h008111,h008112),
       H008102(h008102,dbv0,dbv0),
       H008201(h008201,h008211,h008212),
       H008202(h008202,dbv0,dbv0),
       H008301(h008301,h008311,h008312),
       H008302(h008302,dbv0,dbv0),
       H008401(h008401,h008411,h008412),
       H008402(h008402,dbv0,dbv0),
       H008501(h008501,h008511,h008512),
       H008502(h008502,dbv0,dbv0),
       H008601(h008601,h008611,h008612),
       H008602(h008602,dbv0,dbv0),
       H008701(h008701,h008711,h008712),
       H008702(h008702,dbv0,dbv0),
       H008801(h008801,h008811,h008812),
       H008802(h008802,dbv0,dbv0),
       H008901(h008901,h008911,h008912),
       H008902(h008902,dbv0,dbv0),
       H009001(h009001,h009011,h009012),
       H009002(h009002,dbv0,dbv0);

and    H006111(h006111,h006121,q0061),
       H006112(h006112,h006102,dbv1),
       H006211(h006211,h006221,q0062),
       H006212(h006212,h006202,dbv1),
       H006311(h006311,h006321,q0063),
       H006312(h006312,h006302,dbv1),
       H006411(h006411,h006421,q0064),
       H006412(h006412,h006402,dbv1),
       H006511(h006511,h006521,q0065),
       H006512(h006512,h006502,dbv1),
       H006611(h006611,h006621,q0066),
       H006612(h006612,h006602,dbv1),
       H006711(h006711,h006721,q0067),
       H006712(h006712,h006702,dbv1),
       H006811(h006811,h006821,q0068),
       H006812(h006812,h006802,dbv1),
       H006911(h006911,h006921,q0069),
       H006912(h006912,h006902,dbv1),
       H007011(h007011,h007021,q0070),
       H007012(h007012,h007002,dbv1),
       H007111(h007111,h007121,q0071),
       H007112(h007112,h007102,dbv1),
       H007211(h007211,h007221,q0072),
       H007212(h007212,h007202,dbv1),
       H007311(h007311,h007321,q0073),
       H007312(h007312,h007302,dbv1),
       H007411(h007411,h007421,q0074),
       H007412(h007412,h007402,dbv1),
       H007511(h007511,h007521,q0075),
       H007512(h007512,h007502,dbv1),
       H007611(h007611,h007621,q0076),
       H007612(h007612,h007602,dbv1),
       H007711(h007711,h007721,q0077),
       H007712(h007712,h007702,dbv1),
       H007811(h007811,h007821,q0078),
       H007812(h007812,h007802,dbv1),
       H007911(h007911,h007921,q0079),
       H007912(h007912,h007902,dbv1),
       H008011(h008011,h008021,q0080),
       H008012(h008012,h008002,dbv1),
       H008111(h008111,h008121,q0081),
       H008112(h008112,h008102,dbv0),
       H008211(h008211,h008221,q0082),
       H008212(h008212,h008202,dbv0),
       H008311(h008311,h008321,q0083),
       H008312(h008312,h008302,dbv0),
       H008411(h008411,h008421,q0084),
       H008412(h008412,h008402,dbv0),
       H008511(h008511,h008521,q0085),
       H008512(h008512,h008502,dbv0),
       H008611(h008611,h008621,q0086),
       H008612(h008612,h008602,dbv0),
       H008711(h008711,h008721,q0087),
       H008712(h008712,h008702,dbv0),
       H008811(h008811,h008821,q0088),
       H008812(h008812,h008802,dbv0),
       H008911(h008911,h008921,q0089),
       H008912(h008912,h008902,dbv0),
       H009011(h009011,h009021,q0090),
       H009012(h009012,h009002,dbv0);

not    H006121(h006121,h006102),
       H006221(h006221,h006202),
       H006321(h006321,h006302),
       H006421(h006421,h006402),
       H006521(h006521,h006502),
       H006621(h006621,h006602),
       H006721(h006721,h006702),
       H006821(h006821,h006802),
       H006921(h006921,h006902),
       H007021(h007021,h007002),
       H007121(h007121,h007102),
       H007221(h007221,h007202),
       H007321(h007321,h007302),
       H007421(h007421,h007402),
       H007521(h007521,h007502),
       H007621(h007621,h007602),
       H007721(h007721,h007702),
       H007821(h007821,h007802),
       H007921(h007921,h007902),
       H008021(h008021,h008002),
       H008121(h008121,h008102),
       H008221(h008221,h008202),
       H008321(h008321,h008302),
       H008421(h008421,h008402),
       H008521(h008521,h008502),
       H008621(h008621,h008602),
       H008721(h008721,h008702),
       H008821(h008821,h008802),
       H008921(h008921,h008902),
       H009021(h009021,h009002);

or     O3190(o3190,x0061,x0062,x0063,x0064,x0065,x0066,x0067,x0068,x0069,x0070,x0071,x0072,x0073,x0074,x0075,x0076,x0077,x0078,x0079,x0080,x0081,x0082,x0083,x0084,x0085,x0086,x0087,x0088,x0089,x0090);
not    N3190(n3190,o3190);
//y
not    N0091(n0091,q0091);
xor    X0092(x0092,q0092,q0091),
       X0093(x0093,q0093,a0093),
       X0094(x0094,q0094,a0094),
       X0095(x0095,q0095,a0095),
       X0096(x0096,q0096,a0096),
       X0097(x0097,q0097,a0097),
       X0098(x0098,q0098,a0098),
       X0099(x0099,q0099,a0099),
       X0100(x0100,q0100,a0100),
       X0101(x0101,q0101,a0101),
       X0102(x0102,q0102,a0102),
       X0103(x0103,q0103,a0103),
       X0104(x0104,q0104,a0104),
       X0105(x0105,q0105,a0105),
       X0106(x0106,q0106,a0106),
       X0107(x0107,q0107,a0107),
       X0108(x0108,q0108,a0108),
       X0109(x0109,q0109,a0109),
       X0110(x0110,q0110,a0110),
       X0111(x0111,q0111,a0111),
       X0112(x0112,q0112,a0112),
       X0113(x0113,q0113,a0113),
       X0114(x0114,q0114,a0114),
       X0115(x0115,q0115,a0115),
       X0116(x0116,q0116,a0116),
       X0117(x0117,q0117,a0117),
       X0118(x0118,q0118,a0118),
       X0119(x0119,q0119,a0119),
       X0120(x0120,q0120,a0120);

and    A0093(a0093,q0092,q0091),
       A0094(a0094,a0093,q0093),
       A0095(a0095,a0094,q0094),
       A0096(a0096,a0095,q0095),
       A0097(a0097,a0096,q0096),
       A0098(a0098,a0097,q0097),
       A0099(a0099,a0098,q0098),
       A0100(a0100,a0099,q0099),
       A0101(a0101,a0100,q0100),
       A0102(a0102,a0101,q0101),
       A0103(a0103,a0102,q0102),
       A0104(a0104,a0103,q0103),
       A0105(a0105,a0104,q0104),
       A0106(a0106,a0105,q0105),
       A0107(a0107,a0106,q0106),
       A0108(a0108,a0107,q0107),
       A0109(a0109,a0108,q0108),
       A0110(a0110,a0109,q0109),
       A0111(a0111,a0110,q0110),
       A0112(a0112,a0111,q0111),
       A0113(a0113,a0112,q0112),
       A0114(a0114,a0113,q0113),
       A0115(a0115,a0114,q0114),
       A0116(a0116,a0115,q0115),
       A0117(a0117,a0116,q0116),
       A0118(a0118,a0117,q0117),
       A0119(a0119,a0118,q0118),
       A0120(a0120,a0119,q0119);

xor    X0121(x0121,q0121,q0091),
       X0122(x0122,q0122,q0092),
       X0123(x0123,q0123,q0093),
       X0124(x0124,q0124,q0094),
       X0125(x0125,q0125,q0095),
       X0126(x0126,q0126,q0096),
       X0127(x0127,q0127,q0097),
       X0128(x0128,q0128,q0098),
       X0129(x0129,q0129,q0099),
       X0130(x0130,q0130,q0100),
       X0131(x0131,q0131,q0101),
       X0132(x0132,q0132,q0102),
       X0133(x0133,q0133,q0103),
       X0134(x0134,q0134,q0104),
       X0135(x0135,q0135,q0105),
       X0136(x0136,q0136,q0106),
       X0137(x0137,q0137,q0107),
       X0138(x0138,q0138,q0108),
       X0139(x0139,q0139,q0109),
       X0140(x0140,q0140,q0110),
       X0141(x0141,q0141,q0111),
       X0142(x0142,q0142,q0112),
       X0143(x0143,q0143,q0113),
       X0144(x0144,q0144,q0114),
       X0145(x0145,q0145,q0115),
       X0146(x0146,q0146,q0116),
       X0147(x0147,q0147,q0117),
       X0148(x0148,q0148,q0118),
       X0149(x0149,q0149,q0119),
       X0150(x0150,q0150,q0120);

and    A0121(a0121,n0091,o9150,h0_021,n11_1),
       A0122(a0122,x0092,o9150,h0_021,n11_1),
       A0123(a0123,x0093,o9150,h0_021,n11_1),
       A0124(a0124,x0094,o9150,h0_021,n11_1),
       A0125(a0125,x0095,o9150,h0_021,n11_1),
       A0126(a0126,x0096,o9150,h0_021,n11_1),
       A0127(a0127,x0097,o9150,h0_021,n11_1),
       A0128(a0128,x0098,o9150,h0_021,n11_1),
       A0129(a0129,x0099,o9150,h0_021,n11_1),
       A0130(a0130,x0100,o9150,h0_021,n11_1),
       A0131(a0131,x0101,o9150,h0_021,n11_1),
       A0132(a0132,x0102,o9150,h0_021,n11_1),
       A0133(a0133,x0103,o9150,h0_021,n11_1),
       A0134(a0134,x0104,o9150,h0_021,n11_1),
       A0135(a0135,x0105,o9150,h0_021,n11_1),
       A0136(a0136,x0106,o9150,h0_021,n11_1),
       A0137(a0137,x0107,o9150,h0_021,n11_1),
       A0138(a0138,x0108,o9150,h0_021,n11_1),
       A0139(a0139,x0109,o9150,h0_021,n11_1),
       A0140(a0140,x0110,o9150,h0_021,n11_1),
       A0141(a0141,x0111,o9150,h0_021,n11_1),
       A0142(a0142,x0112,o9150,h0_021,n11_1),
       A0143(a0143,x0113,o9150,h0_021,n11_1),
       A0144(a0144,x0114,o9150,h0_021,n11_1),
       A0145(a0145,x0115,o9150,h0_021,n11_1),
       A0146(a0146,x0116,o9150,h0_021,n11_1),
       A0147(a0147,x0117,o9150,h0_021,n11_1),
       A0148(a0148,x0118,o9150,h0_021,n11_1),
       A0149(a0149,x0119,o9150,h0_021,n11_1),
       A0150(a0150,x0120,o9150,h0_021,n11_1);

or     H012101(h012101,h012111,h012112,q11_1),
       H012102(h012102,h0_002,h0_002,q11_1),
       H012201(h012201,h012211,h012212,q11_1),
       H012202(h012202,h0_002,h0_002,q11_1),
       H012301(h012301,h012311,h012312,q11_1),
       H012302(h012302,h0_002,h0_002,q11_1),
       H012401(h012401,h012411,h012412,q11_1),
       H012402(h012402,h0_002,h0_002,q11_1),
       H012501(h012501,h012511,h012512,q11_1),
       H012502(h012502,h0_002,h0_002,q11_1),
       H012601(h012601,h012611,h012612,q11_1),
       H012602(h012602,h0_002,h0_002,q11_1),
       H012701(h012701,h012711,h012712,q11_1),
       H012702(h012702,h0_002,h0_002,q11_1),
       H012801(h012801,h012811,h012812,q11_1),
       H012802(h012802,h0_002,h0_002,q11_1),
       H012901(h012901,h012911,h012912,q11_1),
       H012902(h012902,h0_002,h0_002,q11_1),
       H013001(h013001,h013011,h013012,q11_1),
       H013002(h013002,h0_002,h0_002,q11_1),
       H013101(h013101,h013111,h013112,q11_1),
       H013102(h013102,h0_002,h0_002,q11_1),
       H013201(h013201,h013211,h013212,q11_1),
       H013202(h013202,h0_002,h0_002,q11_1),
       H013301(h013301,h013311,h013312,q11_1),
       H013302(h013302,h0_002,h0_002,q11_1),
       H013401(h013401,h013411,h013412,q11_1),
       H013402(h013402,h0_002,h0_002,q11_1),
       H013501(h013501,h013511,h013512,q11_1),
       H013502(h013502,h0_002,h0_002,q11_1),
       H013601(h013601,h013611,h013612,q11_1),
       H013602(h013602,h0_002,h0_002,q11_1),
       H013701(h013701,h013711,h013712,q11_1),
       H013702(h013702,h0_002,h0_002,q11_1),
       H013801(h013801,h013811,h013812,q11_1),
       H013802(h013802,h0_002,h0_002,q11_1),
       H013901(h013901,h013911,h013912,q11_1),
       H013902(h013902,h0_002,h0_002,q11_1),
       H014001(h014001,h014011,h014012,q11_1),
       H014002(h014002,h0_002,h0_002,q11_1),
       H014101(h014101,h014111,h014112,q11_1),
       H014102(h014102,h0_002,h0_002,q11_1),
       H014201(h014201,h014211,h014212,q11_1),
       H014202(h014202,h0_002,h0_002,q11_1),
       H014301(h014301,h014311,h014312,q11_1),
       H014302(h014302,h0_002,h0_002,q11_1),
       H014401(h014401,h014411,h014412),
       H014402(h014402,h0_002,h0_002),
       H014501(h014501,h014511,h014512),
       H014502(h014502,h0_002,h0_002),
       H014601(h014601,h014611,h014612),
       H014602(h014602,h0_002,h0_002),
       H014701(h014701,h014711,h014712),
       H014702(h014702,h0_002,h0_002),
       H014801(h014801,h014811,h014812),
       H014802(h014802,h0_002,h0_002),
       H014901(h014901,h014911,h014912),
       H014902(h014902,h0_002,h0_002),
       H015001(h015001,h015011,h015012),
       H015002(h015002,h0_002,h0_002);

and    H012111(h012111,h012121,q0121),
       H012112(h012112,h012102,dbv1),
       H012211(h012211,h012221,q0122),
       H012212(h012212,h012202,dbv1),
       H012311(h012311,h012321,q0123),
       H012312(h012312,h012302,dbv1),
       H012411(h012411,h012421,q0124),
       H012412(h012412,h012402,dbv1),
       H012511(h012511,h012521,q0125),
       H012512(h012512,h012502,dbv1),
       H012611(h012611,h012621,q0126),
       H012612(h012612,h012602,dbv1),
       H012711(h012711,h012721,q0127),
       H012712(h012712,h012702,dbv1),
       H012811(h012811,h012821,q0128),
       H012812(h012812,h012802,dbv1),
       H012911(h012911,h012921,q0129),
       H012912(h012912,h012902,q29_0),
       H013011(h013011,h013021,q0130),
       H013012(h013012,h013002,q30_0),
       H013111(h013111,h013121,q0131),
       H013112(h013112,h013102,q31_0),
       H013211(h013211,h013221,q0132),
       H013212(h013212,h013202,q32_0),
       H013311(h013311,h013321,q0133),
       H013312(h013312,h013302,q33_0),
       H013411(h013411,h013421,q0134),
       H013412(h013412,h013402,q34_0),
       H013511(h013511,h013521,q0135),
       H013512(h013512,h013502,q35_0),
       H013611(h013611,h013621,q0136),
       H013612(h013612,h013602,q36_0),
       H013711(h013711,h013721,q0137),
       H013712(h013712,h013702,q37_0),
       H013811(h013811,h013821,q0138),
       H013812(h013812,h013802,q38_0),
       H013911(h013911,h013921,q0139),
       H013912(h013912,h013902,q39_0),
       H014011(h014011,h014021,q0140),
       H014012(h014012,h014002,q40_0),
       H014111(h014111,h014121,q0141),
       H014112(h014112,h014102,q41_0),
       H014211(h014211,h014221,q0142),
       H014212(h014212,h014202,q42_0),
       H014311(h014311,h014321,q0143),
       H014312(h014312,h014302,q43_0),
       H014411(h014411,h014421,q0144),
       H014412(h014412,h014402,q44_0),
       H014511(h014511,h014521,q0145),
       H014512(h014512,h014502,q45_0),
       H014611(h014611,h014621,q0146),
       H014612(h014612,h014602,q46_0),
       H014711(h014711,h014721,q0147),
       H014712(h014712,h014702,q47_0),
       H014811(h014811,h014821,q0148),
       H014812(h014812,h014802,q48_0),
       H014911(h014911,h014921,q0149),
       H014912(h014912,h014902,q49_0),
       H015011(h015011,h015021,q0150),
       H015012(h015012,h015002,q50_0);

not    H012121(h012121,h012102),
       H012221(h012221,h012202),
       H012321(h012321,h012302),
       H012421(h012421,h012402),
       H012521(h012521,h012502),
       H012621(h012621,h012602),
       H012721(h012721,h012702),
       H012821(h012821,h012802),
       H012921(h012921,h012902),
       H013021(h013021,h013002),
       H013121(h013121,h013102),
       H013221(h013221,h013202),
       H013321(h013321,h013302),
       H013421(h013421,h013402),
       H013521(h013521,h013502),
       H013621(h013621,h013602),
       H013721(h013721,h013702),
       H013821(h013821,h013802),
       H013921(h013921,h013902),
       H014021(h014021,h014002),
       H014121(h014121,h014102),
       H014221(h014221,h014202),
       H014321(h014321,h014302),
       H014421(h014421,h014402),
       H014521(h014521,h014502),
       H014621(h014621,h014602),
       H014721(h014721,h014702),
       H014821(h014821,h014802),
       H014921(h014921,h014902),
       H015021(h015021,h015002);

or     O9150(o9150,x0121,x0122,x0123,x0124,x0125,x0126,x0127,x0128,x0129,x0130,x0131,x0132,x0133,x0134,x0135,x0136,x0137,x0138,x0139,x0140,x0141,x0142,x0143,x0144,x0145,x0146,x0147,x0148,x0149,x0150);
not    N9150(n9150,o9150);
//1
not    N0151(n0151,q0151);
xor    X0152(x0152,q0152,q0151),
       X0153(x0153,q0153,a0153),
       X0154(x0154,q0154,a0154),
       X0155(x0155,q0155,a0155),
       X0156(x0156,q0156,a0156),
       X0157(x0157,q0157,a0157),
       X0158(x0158,q0158,a0158),
       X0159(x0159,q0159,a0159),
       X0160(x0160,q0160,a0160),
       X0161(x0161,q0161,a0161),
       X0162(x0162,q0162,a0162),
       X0163(x0163,q0163,a0163),
       X0164(x0164,q0164,a0164),
       X0165(x0165,q0165,a0165),
       X0166(x0166,q0166,a0166),
       X0167(x0167,q0167,a0167),
       X0168(x0168,q0168,a0168),
       X0169(x0169,q0169,a0169),
       X0170(x0170,q0170,a0170),
       X0171(x0171,q0171,a0171),
       X0172(x0172,q0172,a0172),
       X0173(x0173,q0173,a0173),
       X0174(x0174,q0174,a0174),
       X0175(x0175,q0175,a0175),
       X0176(x0176,q0176,a0176),
       X0177(x0177,q0177,a0177),
       X0178(x0178,q0178,a0178),
       X0179(x0179,q0179,a0179),
       X0180(x0180,q0180,a0180);

and    A0153(a0153,q0152,q0151),
       A0154(a0154,a0153,q0153),
       A0155(a0155,a0154,q0154),
       A0156(a0156,a0155,q0155),
       A0157(a0157,a0156,q0156),
       A0158(a0158,a0157,q0157),
       A0159(a0159,a0158,q0158),
       A0160(a0160,a0159,q0159),
       A0161(a0161,a0160,q0160),
       A0162(a0162,a0161,q0161),
       A0163(a0163,a0162,q0162),
       A0164(a0164,a0163,q0163),
       A0165(a0165,a0164,q0164),
       A0166(a0166,a0165,q0165),
       A0167(a0167,a0166,q0166),
       A0168(a0168,a0167,q0167),
       A0169(a0169,a0168,q0168),
       A0170(a0170,a0169,q0169),
       A0171(a0171,a0170,q0170),
       A0172(a0172,a0171,q0171),
       A0173(a0173,a0172,q0172),
       A0174(a0174,a0173,q0173),
       A0175(a0175,a0174,q0174),
       A0176(a0176,a0175,q0175),
       A0177(a0177,a0176,q0176),
       A0178(a0178,a0177,q0177),
       A0179(a0179,a0178,q0178),
       A0180(a0180,a0179,q0179);

xor    X0181(x0181,q0181,q0151),
       X0182(x0182,q0182,q0152),
       X0183(x0183,q0183,q0153),
       X0184(x0184,q0184,q0154),
       X0185(x0185,q0185,q0155),
       X0186(x0186,q0186,q0156),
       X0187(x0187,q0187,q0157),
       X0188(x0188,q0188,q0158),
       X0189(x0189,q0189,q0159),
       X0190(x0190,q0190,q0160),
       X0191(x0191,q0191,q0161),
       X0192(x0192,q0192,q0162),
       X0193(x0193,q0193,q0163),
       X0194(x0194,q0194,q0164),
       X0195(x0195,q0195,q0165),
       X0196(x0196,q0196,q0166),
       X0197(x0197,q0197,q0167),
       X0198(x0198,q0198,q0168),
       X0199(x0199,q0199,q0169),
       X0200(x0200,q0200,q0170),
       X0201(x0201,q0201,q0171),
       X0202(x0202,q0202,q0172),
       X0203(x0203,q0203,q0173),
       X0204(x0204,q0204,q0174),
       X0205(x0205,q0205,q0175),
       X0206(x0206,q0206,q0176),
       X0207(x0207,q0207,q0177),
       X0208(x0208,q0208,q0178),
       X0209(x0209,q0209,q0179),
       X0210(x0210,q0210,q0180);

and    A0181(a0181,n0151,o5110,xs),
       A0182(a0182,x0152,o5110,xs),
       A0183(a0183,x0153,o5110,xs),
       A0184(a0184,x0154,o5110,xs),
       A0185(a0185,x0155,o5110,xs),
       A0186(a0186,x0156,o5110,xs),
       A0187(a0187,x0157,o5110,xs),
       A0188(a0188,x0158,o5110,xs),
       A0189(a0189,x0159,o5110,xs),
       A0190(a0190,x0160,o5110,xs),
       A0191(a0191,x0161,o5110,xs),
       A0192(a0192,x0162,o5110,xs),
       A0193(a0193,x0163,o5110,xs),
       A0194(a0194,x0164,o5110,xs),
       A0195(a0195,x0165,o5110,xs),
       A0196(a0196,x0166,o5110,xs),
       A0197(a0197,x0167,o5110,xs),
       A0198(a0198,x0168,o5110,xs),
       A0199(a0199,x0169,o5110,xs),
       A0200(a0200,x0170,o5110,xs),
       A0201(a0201,x0171,o5110,xs),
       A0202(a0202,x0172,o5110,xs),
       A0203(a0203,x0173,o5110,xs),
       A0204(a0204,x0174,o5110,xs),
       A0205(a0205,x0175,o5110,xs),
       A0206(a0206,x0176,o5110,xs),
       A0207(a0207,x0177,o5110,xs),
       A0208(a0208,x0178,o5110,xs),
       A0209(a0209,x0179,o5110,xs),
       A0210(a0210,x0180,o5110,xs);

or     H018101(h018101,h018111,h018112),
       H018102(h018102,dbv0,dbv0),
       H018201(h018201,h018211,h018212),
       H018202(h018202,dbv0,dbv0),
       H018301(h018301,h018311,h018312),
       H018302(h018302,dbv0,dbv0),
       H018401(h018401,h018411,h018412),
       H018402(h018402,dbv0,dbv0),
       H018501(h018501,h018511,h018512),
       H018502(h018502,dbv0,dbv0),
       H018601(h018601,h018611,h018612),
       H018602(h018602,dbv0,dbv0),
       H018701(h018701,h018711,h018712),
       H018702(h018702,dbv0,dbv0),
       H018801(h018801,h018811,h018812),
       H018802(h018802,dbv0,dbv0),
       H018901(h018901,h018911,h018912),
       H018902(h018902,dbv0,dbv0),
       H019001(h019001,h019011,h019012),
       H019002(h019002,dbv0,dbv0),
       H019101(h019101,h019111,h019112),
       H019102(h019102,dbv0,dbv0),
       H019201(h019201,h019211,h019212),
       H019202(h019202,dbv0,dbv0),
       H019301(h019301,h019311,h019312),
       H019302(h019302,dbv0,dbv0),
       H019401(h019401,h019411,h019412),
       H019402(h019402,dbv0,dbv0),
       H019501(h019501,h019511,h019512),
       H019502(h019502,dbv0,dbv0),
       H019601(h019601,h019611,h019612),
       H019602(h019602,dbv0,dbv0),
       H019701(h019701,h019711,h019712),
       H019702(h019702,dbv0,dbv0),
       H019801(h019801,h019811,h019812),
       H019802(h019802,dbv0,dbv0),
       H019901(h019901,h019911,h019912),
       H019902(h019902,dbv0,dbv0),
       H020001(h020001,h020011,h020012),
       H020002(h020002,dbv0,dbv0),
       H020101(h020101,h020111,h020112),
       H020102(h020102,dbv0,dbv0),
       H020201(h020201,h020211,h020212),
       H020202(h020202,dbv0,dbv0),
       H020301(h020301,h020311,h020312),
       H020302(h020302,dbv0,dbv0),
       H020401(h020401,h020411,h020412),
       H020402(h020402,dbv0,dbv0),
       H020501(h020501,h020511,h020512),
       H020502(h020502,dbv0,dbv0),
       H020601(h020601,h020611,h020612),
       H020602(h020602,dbv0,dbv0),
       H020701(h020701,h020711,h020712),
       H020702(h020702,dbv0,dbv0),
       H020801(h020801,h020811,h020812),
       H020802(h020802,dbv0,dbv0),
       H020901(h020901,h020911,h020912),
       H020902(h020902,dbv0,dbv0),
       H021001(h021001,h021011,h021012),
       H021002(h021002,dbv0,dbv0);

and    H018111(h018111,h018121,q0181),
       H018112(h018112,h018102,q0181),
       H018211(h018211,h018221,q0182),
       H018212(h018212,h018202,q0182),
       H018311(h018311,h018321,q0183),
       H018312(h018312,h018302,q0183),
       H018411(h018411,h018421,q0184),
       H018412(h018412,h018402,q0184),
       H018511(h018511,h018521,q0185),
       H018512(h018512,h018502,q0185),
       H018611(h018611,h018621,q0186),
       H018612(h018612,h018602,q0186),
       H018711(h018711,h018721,q0187),
       H018712(h018712,h018702,q0187),
       H018811(h018811,h018821,q0188),
       H018812(h018812,h018802,q0188),
       H018911(h018911,h018921,q0189),
       H018912(h018912,h018902,q0189),
       H019011(h019011,h019021,q0190),
       H019012(h019012,h019002,q0190),
       H019111(h019111,h019121,q0191),
       H019112(h019112,h019102,q0191),
       H019211(h019211,h019221,q0192),
       H019212(h019212,h019202,q0192),
       H019311(h019311,h019321,q0193),
       H019312(h019312,h019302,q0193),
       H019411(h019411,h019421,q0194),
       H019412(h019412,h019402,q0194),
       H019511(h019511,h019521,q0195),
       H019512(h019512,h019502,q0195),
       H019611(h019611,h019621,q0196),
       H019612(h019612,h019602,q0196),
       H019711(h019711,h019721,q0197),
       H019712(h019712,h019702,q0197),
       H019811(h019811,h019821,q0198),
       H019812(h019812,h019802,q0198),
       H019911(h019911,h019921,q0199),
       H019912(h019912,h019902,q0199),
       H020011(h020011,h020021,q0200),
       H020012(h020012,h020002,q0200),
       H020111(h020111,h020121,q0201),
       H020112(h020112,h020102,q0201),
       H020211(h020211,h020221,q0202),
       H020212(h020212,h020202,q0202),
       H020311(h020311,h020321,q0203),
       H020312(h020312,h020302,q0203),
       H020411(h020411,h020421,q0204),
       H020412(h020412,h020402,q0204),
       H020511(h020511,h020521,q0205),
       H020512(h020512,h020502,q0205),
       H020611(h020611,h020621,q0206),
       H020612(h020612,h020602,q0206),
       H020711(h020711,h020721,q0207),
       H020712(h020712,h020702,q0207),
       H020811(h020811,h020821,q0208),
       H020812(h020812,h020802,q0208),
       H020911(h020911,h020921,q0209),
       H020912(h020912,h020902,q0209),
       H021011(h021011,h021021,q0210),
       H021012(h021012,h021002,q0210);

not    H018121(h018121,h018102),
       H018221(h018221,h018202),
       H018321(h018321,h018302),
       H018421(h018421,h018402),
       H018521(h018521,h018502),
       H018621(h018621,h018602),
       H018721(h018721,h018702),
       H018821(h018821,h018802),
       H018921(h018921,h018902),
       H019021(h019021,h019002),
       H019121(h019121,h019102),
       H019221(h019221,h019202),
       H019321(h019321,h019302),
       H019421(h019421,h019402),
       H019521(h019521,h019502),
       H019621(h019621,h019602),
       H019721(h019721,h019702),
       H019821(h019821,h019802),
       H019921(h019921,h019902),
       H020021(h020021,h020002),
       H020121(h020121,h020102),
       H020221(h020221,h020202),
       H020321(h020321,h020302),
       H020421(h020421,h020402),
       H020521(h020521,h020502),
       H020621(h020621,h020602),
       H020721(h020721,h020702),
       H020821(h020821,h020802),
       H020921(h020921,h020902),
       H021021(h021021,h021002);

or     O5110(o5110,x0181,x0182,x0183,x0184,x0185,x0186,x0187,x0188,x0189,x0190,x0191,x0192,x0193,x0194,x0195,x0196,x0197,x0198,x0199,x0200,x0201,x0202,x0203,x0204,x0205,x0206,x0207,x0208,x0209,x0210);
not    N5110(n5110,o5110);
//2
not    N0211(n0211,q0211);
xor    X0212(x0212,q0212,q0211),
       X0213(x0213,q0213,a0213),
       X0214(x0214,q0214,a0214),
       X0215(x0215,q0215,a0215),
       X0216(x0216,q0216,a0216),
       X0217(x0217,q0217,a0217),
       X0218(x0218,q0218,a0218),
       X0219(x0219,q0219,a0219),
       X0220(x0220,q0220,a0220),
       X0221(x0221,q0221,a0221),
       X0222(x0222,q0222,a0222),
       X0223(x0223,q0223,a0223),
       X0224(x0224,q0224,a0224),
       X0225(x0225,q0225,a0225),
       X0226(x0226,q0226,a0226),
       X0227(x0227,q0227,a0227),
       X0228(x0228,q0228,a0228),
       X0229(x0229,q0229,a0229),
       X0230(x0230,q0230,a0230),
       X0231(x0231,q0231,a0231),
       X0232(x0232,q0232,a0232),
       X0233(x0233,q0233,a0233),
       X0234(x0234,q0234,a0234),
       X0235(x0235,q0235,a0235),
       X0236(x0236,q0236,a0236),
       X0237(x0237,q0237,a0237),
       X0238(x0238,q0238,a0238),
       X0239(x0239,q0239,a0239),
       X0240(x0240,q0240,a0240);

and    A0213(a0213,q0212,q0211),
       A0214(a0214,a0213,q0213),
       A0215(a0215,a0214,q0214),
       A0216(a0216,a0215,q0215),
       A0217(a0217,a0216,q0216),
       A0218(a0218,a0217,q0217),
       A0219(a0219,a0218,q0218),
       A0220(a0220,a0219,q0219),
       A0221(a0221,a0220,q0220),
       A0222(a0222,a0221,q0221),
       A0223(a0223,a0222,q0222),
       A0224(a0224,a0223,q0223),
       A0225(a0225,a0224,q0224),
       A0226(a0226,a0225,q0225),
       A0227(a0227,a0226,q0226),
       A0228(a0228,a0227,q0227),
       A0229(a0229,a0228,q0228),
       A0230(a0230,a0229,q0229),
       A0231(a0231,a0230,q0230),
       A0232(a0232,a0231,q0231),
       A0233(a0233,a0232,q0232),
       A0234(a0234,a0233,q0233),
       A0235(a0235,a0234,q0234),
       A0236(a0236,a0235,q0235),
       A0237(a0237,a0236,q0236),
       A0238(a0238,a0237,q0237),
       A0239(a0239,a0238,q0238),
       A0240(a0240,a0239,q0239);

xor    X0241(x0241,q0241,q0211),
       X0242(x0242,q0242,q0212),
       X0243(x0243,q0243,q0213),
       X0244(x0244,q0244,q0214),
       X0245(x0245,q0245,q0215),
       X0246(x0246,q0246,q0216),
       X0247(x0247,q0247,q0217),
       X0248(x0248,q0248,q0218),
       X0249(x0249,q0249,q0219),
       X0250(x0250,q0250,q0220),
       X0251(x0251,q0251,q0221),
       X0252(x0252,q0252,q0222),
       X0253(x0253,q0253,q0223),
       X0254(x0254,q0254,q0224),
       X0255(x0255,q0255,q0225),
       X0256(x0256,q0256,q0226),
       X0257(x0257,q0257,q0227),
       X0258(x0258,q0258,q0228),
       X0259(x0259,q0259,q0229),
       X0260(x0260,q0260,q0230),
       X0261(x0261,q0261,q0231),
       X0262(x0262,q0262,q0232),
       X0263(x0263,q0263,q0233),
       X0264(x0264,q0264,q0234),
       X0265(x0265,q0265,q0235),
       X0266(x0266,q0266,q0236),
       X0267(x0267,q0267,q0237),
       X0268(x0268,q0268,q0238),
       X0269(x0269,q0269,q0239),
       X0270(x0270,q0270,q0240);

and    A0241(a0241,n0211,o1170,xk),
       A0242(a0242,x0212,o1170,xk),
       A0243(a0243,x0213,o1170,xk),
       A0244(a0244,x0214,o1170,xk),
       A0245(a0245,x0215,o1170,xk),
       A0246(a0246,x0216,o1170,xk),
       A0247(a0247,x0217,o1170,xk),
       A0248(a0248,x0218,o1170,xk),
       A0249(a0249,x0219,o1170,xk),
       A0250(a0250,x0220,o1170,xk),
       A0251(a0251,x0221,o1170,xk),
       A0252(a0252,x0222,o1170,xk),
       A0253(a0253,x0223,o1170,xk),
       A0254(a0254,x0224,o1170,xk),
       A0255(a0255,x0225,o1170,xk),
       A0256(a0256,x0226,o1170,xk),
       A0257(a0257,x0227,o1170,xk),
       A0258(a0258,x0228,o1170,xk),
       A0259(a0259,x0229,o1170,xk),
       A0260(a0260,x0230,o1170,xk),
       A0261(a0261,x0231,o1170,xk),
       A0262(a0262,x0232,o1170,xk),
       A0263(a0263,x0233,o1170,xk),
       A0264(a0264,x0234,o1170,xk),
       A0265(a0265,x0235,o1170,xk),
       A0266(a0266,x0236,o1170,xk),
       A0267(a0267,x0237,o1170,xk),
       A0268(a0268,x0238,o1170,xk),
       A0269(a0269,x0239,o1170,xk),
       A0270(a0270,x0240,o1170,xk);

or     H024101(h024101,h024111,h024112),
       H024102(h024102,dbv0,dbv0),
       H024201(h024201,h024211,h024212),
       H024202(h024202,dbv0,dbv0),
       H024301(h024301,h024311,h024312),
       H024302(h024302,dbv0,dbv0),
       H024401(h024401,h024411,h024412),
       H024402(h024402,dbv0,dbv0),
       H024501(h024501,h024511,h024512),
       H024502(h024502,dbv0,dbv0),
       H024601(h024601,h024611,h024612),
       H024602(h024602,dbv0,dbv0),
       H024701(h024701,h024711,h024712),
       H024702(h024702,dbv0,dbv0),
       H024801(h024801,h024811,h024812),
       H024802(h024802,dbv0,dbv0),
       H024901(h024901,h024911,h024912),
       H024902(h024902,dbv0,dbv0),
       H025001(h025001,h025011,h025012),
       H025002(h025002,dbv0,dbv0),
       H025101(h025101,h025111,h025112),
       H025102(h025102,dbv0,dbv0),
       H025201(h025201,h025211,h025212),
       H025202(h025202,dbv0,dbv0),
       H025301(h025301,h025311,h025312),
       H025302(h025302,dbv0,dbv0),
       H025401(h025401,h025411,h025412),
       H025402(h025402,dbv0,dbv0),
       H025501(h025501,h025511,h025512),
       H025502(h025502,dbv0,dbv0),
       H025601(h025601,h025611,h025612),
       H025602(h025602,dbv0,dbv0),
       H025701(h025701,h025711,h025712),
       H025702(h025702,dbv0,dbv0),
       H025801(h025801,h025811,h025812),
       H025802(h025802,dbv0,dbv0),
       H025901(h025901,h025911,h025912),
       H025902(h025902,dbv0,dbv0),
       H026001(h026001,h026011,h026012),
       H026002(h026002,dbv0,dbv0),
       H026101(h026101,h026111,h026112),
       H026102(h026102,dbv0,dbv0),
       H026201(h026201,h026211,h026212),
       H026202(h026202,dbv0,dbv0),
       H026301(h026301,h026311,h026312),
       H026302(h026302,dbv0,dbv0),
       H026401(h026401,h026411,h026412),
       H026402(h026402,dbv0,dbv0),
       H026501(h026501,h026511,h026512),
       H026502(h026502,dbv0,dbv0),
       H026601(h026601,h026611,h026612),
       H026602(h026602,dbv0,dbv0),
       H026701(h026701,h026711,h026712),
       H026702(h026702,dbv0,dbv0),
       H026801(h026801,h026811,h026812),
       H026802(h026802,dbv0,dbv0),
       H026901(h026901,h026911,h026912),
       H026902(h026902,dbv0,dbv0),
       H027001(h027001,h027011,h027012),
       H027002(h027002,dbv0,dbv0);

and    H024111(h024111,h024121,q0241),
       H024112(h024112,h024102,q0241),
       H024211(h024211,h024221,q0242),
       H024212(h024212,h024202,q0242),
       H024311(h024311,h024321,q0243),
       H024312(h024312,h024302,q0243),
       H024411(h024411,h024421,q0244),
       H024412(h024412,h024402,q0244),
       H024511(h024511,h024521,q0245),
       H024512(h024512,h024502,q0245),
       H024611(h024611,h024621,q0246),
       H024612(h024612,h024602,q0246),
       H024711(h024711,h024721,q0247),
       H024712(h024712,h024702,q0247),
       H024811(h024811,h024821,q0248),
       H024812(h024812,h024802,q0248),
       H024911(h024911,h024921,q0249),
       H024912(h024912,h024902,q0249),
       H025011(h025011,h025021,q0250),
       H025012(h025012,h025002,q0250),
       H025111(h025111,h025121,q0251),
       H025112(h025112,h025102,q0251),
       H025211(h025211,h025221,q0252),
       H025212(h025212,h025202,q0252),
       H025311(h025311,h025321,q0253),
       H025312(h025312,h025302,q0253),
       H025411(h025411,h025421,q0254),
       H025412(h025412,h025402,q0254),
       H025511(h025511,h025521,q0255),
       H025512(h025512,h025502,q0255),
       H025611(h025611,h025621,q0256),
       H025612(h025612,h025602,q0256),
       H025711(h025711,h025721,q0257),
       H025712(h025712,h025702,q0257),
       H025811(h025811,h025821,q0258),
       H025812(h025812,h025802,q0258),
       H025911(h025911,h025921,q0259),
       H025912(h025912,h025902,q0259),
       H026011(h026011,h026021,q0260),
       H026012(h026012,h026002,q0260),
       H026111(h026111,h026121,q0261),
       H026112(h026112,h026102,q0261),
       H026211(h026211,h026221,q0262),
       H026212(h026212,h026202,q0262),
       H026311(h026311,h026321,q0263),
       H026312(h026312,h026302,q0263),
       H026411(h026411,h026421,q0264),
       H026412(h026412,h026402,q0264),
       H026511(h026511,h026521,q0265),
       H026512(h026512,h026502,q0265),
       H026611(h026611,h026621,q0266),
       H026612(h026612,h026602,q0266),
       H026711(h026711,h026721,q0267),
       H026712(h026712,h026702,q0267),
       H026811(h026811,h026821,q0268),
       H026812(h026812,h026802,q0268),
       H026911(h026911,h026921,q0269),
       H026912(h026912,h026902,q0269),
       H027011(h027011,h027021,q0270),
       H027012(h027012,h027002,q0270);

not    H024121(h024121,h024102),
       H024221(h024221,h024202),
       H024321(h024321,h024302),
       H024421(h024421,h024402),
       H024521(h024521,h024502),
       H024621(h024621,h024602),
       H024721(h024721,h024702),
       H024821(h024821,h024802),
       H024921(h024921,h024902),
       H025021(h025021,h025002),
       H025121(h025121,h025102),
       H025221(h025221,h025202),
       H025321(h025321,h025302),
       H025421(h025421,h025402),
       H025521(h025521,h025502),
       H025621(h025621,h025602),
       H025721(h025721,h025702),
       H025821(h025821,h025802),
       H025921(h025921,h025902),
       H026021(h026021,h026002),
       H026121(h026121,h026102),
       H026221(h026221,h026202),
       H026321(h026321,h026302),
       H026421(h026421,h026402),
       H026521(h026521,h026502),
       H026621(h026621,h026602),
       H026721(h026721,h026702),
       H026821(h026821,h026802),
       H026921(h026921,h026902),
       H027021(h027021,h027002);

or     O1170(o1170,x0241,x0242,x0243,x0244,x0245,x0246,x0247,x0248,x0249,x0250,x0251,x0252,x0253,x0254,x0255,x0256,x0257,x0258,x0259,x0260,x0261,x0262,x0263,x0264,x0265,x0266,x0267,x0268,x0269,x0270);
not    N1170(n1170,o1170);
//s
not    N0271(n0271,q0271);
xor    X0272(x0272,q0272,q0271),
       X0273(x0273,q0273,a0273),
       X0274(x0274,q0274,a0274),
       X0275(x0275,q0275,a0275),
       X0276(x0276,q0276,a0276),
       X0277(x0277,q0277,a0277),
       X0278(x0278,q0278,a0278),
       X0279(x0279,q0279,a0279),
       X0280(x0280,q0280,a0280),
       X0281(x0281,q0281,a0281),
       X0282(x0282,q0282,a0282),
       X0283(x0283,q0283,a0283),
       X0284(x0284,q0284,a0284),
       X0285(x0285,q0285,a0285),
       X0286(x0286,q0286,a0286),
       X0287(x0287,q0287,a0287),
       X0288(x0288,q0288,a0288),
       X0289(x0289,q0289,a0289),
       X0290(x0290,q0290,a0290),
       X0291(x0291,q0291,a0291),
       X0292(x0292,q0292,a0292),
       X0293(x0293,q0293,a0293),
       X0294(x0294,q0294,a0294),
       X0295(x0295,q0295,a0295),
       X0296(x0296,q0296,a0296),
       X0297(x0297,q0297,a0297),
       X0298(x0298,q0298,a0298),
       X0299(x0299,q0299,a0299),
       X0300(x0300,q0300,a0300);

and    A0273(a0273,q0272,q0271),
       A0274(a0274,a0273,q0273),
       A0275(a0275,a0274,q0274),
       A0276(a0276,a0275,q0275),
       A0277(a0277,a0276,q0276),
       A0278(a0278,a0277,q0277),
       A0279(a0279,a0278,q0278),
       A0280(a0280,a0279,q0279),
       A0281(a0281,a0280,q0280),
       A0282(a0282,a0281,q0281),
       A0283(a0283,a0282,q0282),
       A0284(a0284,a0283,q0283),
       A0285(a0285,a0284,q0284),
       A0286(a0286,a0285,q0285),
       A0287(a0287,a0286,q0286),
       A0288(a0288,a0287,q0287),
       A0289(a0289,a0288,q0288),
       A0290(a0290,a0289,q0289),
       A0291(a0291,a0290,q0290),
       A0292(a0292,a0291,q0291),
       A0293(a0293,a0292,q0292),
       A0294(a0294,a0293,q0293),
       A0295(a0295,a0294,q0294),
       A0296(a0296,a0295,q0295),
       A0297(a0297,a0296,q0296),
       A0298(a0298,a0297,q0297),
       A0299(a0299,a0298,q0298),
       A0300(a0300,a0299,q0299);

xor    X0301(x0301,q0301,q0271),
       X0302(x0302,q0302,q0272),
       X0303(x0303,q0303,q0273),
       X0304(x0304,q0304,q0274),
       X0305(x0305,q0305,q0275),
       X0306(x0306,q0306,q0276),
       X0307(x0307,q0307,q0277),
       X0308(x0308,q0308,q0278),
       X0309(x0309,q0309,q0279),
       X0310(x0310,q0310,q0280),
       X0311(x0311,q0311,q0281),
       X0312(x0312,q0312,q0282),
       X0313(x0313,q0313,q0283),
       X0314(x0314,q0314,q0284),
       X0315(x0315,q0315,q0285),
       X0316(x0316,q0316,q0286),
       X0317(x0317,q0317,q0287),
       X0318(x0318,q0318,q0288),
       X0319(x0319,q0319,q0289),
       X0320(x0320,q0320,q0290),
       X0321(x0321,q0321,q0291),
       X0322(x0322,q0322,q0292),
       X0323(x0323,q0323,q0293),
       X0324(x0324,q0324,q0294),
       X0325(x0325,q0325,q0295),
       X0326(x0326,q0326,q0296),
       X0327(x0327,q0327,q0297),
       X0328(x0328,q0328,q0298),
       X0329(x0329,q0329,q0299),
       X0330(x0330,q0330,q0300);

and    A0301(a0301,n0271,o7130,qs_1),
       A0302(a0302,x0272,o7130,qs_1),
       A0303(a0303,x0273,o7130,qs_1),
       A0304(a0304,x0274,o7130,qs_1),
       A0305(a0305,x0275,o7130,qs_1),
       A0306(a0306,x0276,o7130,qs_1),
       A0307(a0307,x0277,o7130,qs_1),
       A0308(a0308,x0278,o7130,qs_1),
       A0309(a0309,x0279,o7130,qs_1),
       A0310(a0310,x0280,o7130,qs_1),
       A0311(a0311,x0281,o7130,qs_1),
       A0312(a0312,x0282,o7130,qs_1),
       A0313(a0313,x0283,o7130,qs_1),
       A0314(a0314,x0284,o7130,qs_1),
       A0315(a0315,x0285,o7130,qs_1),
       A0316(a0316,x0286,o7130,qs_1),
       A0317(a0317,x0287,o7130,qs_1),
       A0318(a0318,x0288,o7130,qs_1),
       A0319(a0319,x0289,o7130,qs_1),
       A0320(a0320,x0290,o7130,qs_1),
       A0321(a0321,x0291,o7130,qs_1),
       A0322(a0322,x0292,o7130,qs_1),
       A0323(a0323,x0293,o7130,qs_1),
       A0324(a0324,x0294,o7130,qs_1),
       A0325(a0325,x0295,o7130,qs_1),
       A0326(a0326,x0296,o7130,qs_1),
       A0327(a0327,x0297,o7130,qs_1),
       A0328(a0328,x0298,o7130,qs_1),
       A0329(a0329,x0299,o7130,qs_1),
       A0330(a0330,x0300,o7130,qs_1);

or     H030101(h030101,h030111,h030112),
       H030102(h030102,dbv0,dbv0),
       H030201(h030201,h030211,h030212),
       H030202(h030202,dbv0,dbv0),
       H030301(h030301,h030311,h030312),
       H030302(h030302,dbv0,dbv0),
       H030401(h030401,h030411,h030412),
       H030402(h030402,dbv0,dbv0),
       H030501(h030501,h030511,h030512),
       H030502(h030502,dbv0,dbv0),
       H030601(h030601,h030611,h030612),
       H030602(h030602,dbv0,dbv0),
       H030701(h030701,h030711,h030712),
       H030702(h030702,dbv0,dbv0),
       H030801(h030801,h030811,h030812),
       H030802(h030802,dbv0,dbv0),
       H030901(h030901,h030911,h030912),
       H030902(h030902,dbv0,dbv0),
       H031001(h031001,h031011,h031012),
       H031002(h031002,dbv0,dbv0),
       H031101(h031101,h031111,h031112),
       H031102(h031102,dbv0,dbv0),
       H031201(h031201,h031211,h031212),
       H031202(h031202,dbv0,dbv0),
       H031301(h031301,h031311,h031312),
       H031302(h031302,dbv0,dbv0),
       H031401(h031401,h031411,h031412),
       H031402(h031402,dbv0,dbv0),
       H031501(h031501,h031511,h031512),
       H031502(h031502,dbv0,dbv0),
       H031601(h031601,h031611,h031612),
       H031602(h031602,dbv0,dbv0),
       H031701(h031701,h031711,h031712),
       H031702(h031702,dbv0,dbv0),
       H031801(h031801,h031811,h031812),
       H031802(h031802,dbv0,dbv0),
       H031901(h031901,h031911,h031912),
       H031902(h031902,dbv0,dbv0),
       H032001(h032001,h032011,h032012),
       H032002(h032002,dbv0,dbv0),
       H032101(h032101,h032111,h032112),
       H032102(h032102,dbv0,dbv0),
       H032201(h032201,h032211,h032212),
       H032202(h032202,dbv0,dbv0),
       H032301(h032301,h032311,h032312),
       H032302(h032302,dbv0,dbv0),
       H032401(h032401,h032411,h032412),
       H032402(h032402,dbv0,dbv0),
       H032501(h032501,h032511,h032512),
       H032502(h032502,dbv0,dbv0),
       H032601(h032601,h032611,h032612),
       H032602(h032602,dbv0,dbv0),
       H032701(h032701,h032711,h032712),
       H032702(h032702,dbv0,dbv0),
       H032801(h032801,h032811,h032812),
       H032802(h032802,dbv0,dbv0),
       H032901(h032901,h032911,h032912),
       H032902(h032902,dbv0,dbv0),
       H033001(h033001,h033011,h033012),
       H033002(h033002,dbv0,dbv0);

and    H030111(h030111,h030121,q0301),
       H030112(h030112,h030102,q0301),
       H030211(h030211,h030221,q0302),
       H030212(h030212,h030202,q0302),
       H030311(h030311,h030321,q0303),
       H030312(h030312,h030302,q0303),
       H030411(h030411,h030421,q0304),
       H030412(h030412,h030402,q0304),
       H030511(h030511,h030521,q0305),
       H030512(h030512,h030502,q0305),
       H030611(h030611,h030621,q0306),
       H030612(h030612,h030602,q0306),
       H030711(h030711,h030721,q0307),
       H030712(h030712,h030702,q0307),
       H030811(h030811,h030821,q0308),
       H030812(h030812,h030802,q0308),
       H030911(h030911,h030921,q0309),
       H030912(h030912,h030902,q0309),
       H031011(h031011,h031021,q0310),
       H031012(h031012,h031002,q0310),
       H031111(h031111,h031121,q0311),
       H031112(h031112,h031102,q0311),
       H031211(h031211,h031221,q0312),
       H031212(h031212,h031202,q0312),
       H031311(h031311,h031321,q0313),
       H031312(h031312,h031302,q0313),
       H031411(h031411,h031421,q0314),
       H031412(h031412,h031402,q0314),
       H031511(h031511,h031521,q0315),
       H031512(h031512,h031502,q0315),
       H031611(h031611,h031621,q0316),
       H031612(h031612,h031602,q0316),
       H031711(h031711,h031721,q0317),
       H031712(h031712,h031702,q0317),
       H031811(h031811,h031821,q0318),
       H031812(h031812,h031802,q0318),
       H031911(h031911,h031921,q0319),
       H031912(h031912,h031902,q0319),
       H032011(h032011,h032021,q0320),
       H032012(h032012,h032002,q0320),
       H032111(h032111,h032121,q0321),
       H032112(h032112,h032102,q0321),
       H032211(h032211,h032221,q0322),
       H032212(h032212,h032202,q0322),
       H032311(h032311,h032321,q0323),
       H032312(h032312,h032302,q0323),
       H032411(h032411,h032421,q0324),
       H032412(h032412,h032402,q0324),
       H032511(h032511,h032521,q0325),
       H032512(h032512,h032502,q0325),
       H032611(h032611,h032621,q0326),
       H032612(h032612,h032602,q0326),
       H032711(h032711,h032721,q0327),
       H032712(h032712,h032702,q0327),
       H032811(h032811,h032821,q0328),
       H032812(h032812,h032802,q0328),
       H032911(h032911,h032921,q0329),
       H032912(h032912,h032902,q0329),
       H033011(h033011,h033021,q0330),
       H033012(h033012,h033002,q0330);

not    H030121(h030121,h030102),
       H030221(h030221,h030202),
       H030321(h030321,h030302),
       H030421(h030421,h030402),
       H030521(h030521,h030502),
       H030621(h030621,h030602),
       H030721(h030721,h030702),
       H030821(h030821,h030802),
       H030921(h030921,h030902),
       H031021(h031021,h031002),
       H031121(h031121,h031102),
       H031221(h031221,h031202),
       H031321(h031321,h031302),
       H031421(h031421,h031402),
       H031521(h031521,h031502),
       H031621(h031621,h031602),
       H031721(h031721,h031702),
       H031821(h031821,h031802),
       H031921(h031921,h031902),
       H032021(h032021,h032002),
       H032121(h032121,h032102),
       H032221(h032221,h032202),
       H032321(h032321,h032302),
       H032421(h032421,h032402),
       H032521(h032521,h032502),
       H032621(h032621,h032602),
       H032721(h032721,h032702),
       H032821(h032821,h032802),
       H032921(h032921,h032902),
       H033021(h033021,h033002);

or     O7130(o7130,x0301,x0302,x0303,x0304,x0305,x0306,x0307,x0308,x0309,x0310,x0311,x0312,x0313,x0314,x0315,x0316,x0317,x0318,x0319,x0320,x0321,x0322,x0323,x0324,x0325,x0326,x0327,x0328,x0329,x0330);
not    N7130(n7130,o7130);
//so
not    N0331(n0331,q0331);
xor    X0332(x0332,q0332,q0331),
       X0333(x0333,q0333,a0333),
       X0334(x0334,q0334,a0334),
       X0335(x0335,q0335,a0335),
       X0336(x0336,q0336,a0336),
       X0337(x0337,q0337,a0337),
       X0338(x0338,q0338,a0338),
       X0339(x0339,q0339,a0339),
       X0340(x0340,q0340,a0340),
       X0341(x0341,q0341,a0341),
       X0342(x0342,q0342,a0342),
       X0343(x0343,q0343,a0343),
       X0344(x0344,q0344,a0344),
       X0345(x0345,q0345,a0345),
       X0346(x0346,q0346,a0346),
       X0347(x0347,q0347,a0347),
       X0348(x0348,q0348,a0348),
       X0349(x0349,q0349,a0349),
       X0350(x0350,q0350,a0350),
       X0351(x0351,q0351,a0351),
       X0352(x0352,q0352,a0352),
       X0353(x0353,q0353,a0353),
       X0354(x0354,q0354,a0354),
       X0355(x0355,q0355,a0355),
       X0356(x0356,q0356,a0356),
       X0357(x0357,q0357,a0357),
       X0358(x0358,q0358,a0358),
       X0359(x0359,q0359,a0359),
       X0360(x0360,q0360,a0360);

and    A0333(a0333,q0332,q0331),
       A0334(a0334,a0333,q0333),
       A0335(a0335,a0334,q0334),
       A0336(a0336,a0335,q0335),
       A0337(a0337,a0336,q0336),
       A0338(a0338,a0337,q0337),
       A0339(a0339,a0338,q0338),
       A0340(a0340,a0339,q0339),
       A0341(a0341,a0340,q0340),
       A0342(a0342,a0341,q0341),
       A0343(a0343,a0342,q0342),
       A0344(a0344,a0343,q0343),
       A0345(a0345,a0344,q0344),
       A0346(a0346,a0345,q0345),
       A0347(a0347,a0346,q0346),
       A0348(a0348,a0347,q0347),
       A0349(a0349,a0348,q0348),
       A0350(a0350,a0349,q0349),
       A0351(a0351,a0350,q0350),
       A0352(a0352,a0351,q0351),
       A0353(a0353,a0352,q0352),
       A0354(a0354,a0353,q0353),
       A0355(a0355,a0354,q0354),
       A0356(a0356,a0355,q0355),
       A0357(a0357,a0356,q0356),
       A0358(a0358,a0357,q0357),
       A0359(a0359,a0358,q0358),
       A0360(a0360,a0359,q0359);

xor    X0361(x0361,q0361,q0331),
       X0362(x0362,q0362,q0332),
       X0363(x0363,q0363,q0333),
       X0364(x0364,q0364,q0334),
       X0365(x0365,q0365,q0335),
       X0366(x0366,q0366,q0336),
       X0367(x0367,q0367,q0337),
       X0368(x0368,q0368,q0338),
       X0369(x0369,q0369,q0339),
       X0370(x0370,q0370,q0340),
       X0371(x0371,q0371,q0341),
       X0372(x0372,q0372,q0342),
       X0373(x0373,q0373,q0343),
       X0374(x0374,q0374,q0344),
       X0375(x0375,q0375,q0345),
       X0376(x0376,q0376,q0346),
       X0377(x0377,q0377,q0347),
       X0378(x0378,q0378,q0348),
       X0379(x0379,q0379,q0349),
       X0380(x0380,q0380,q0350),
       X0381(x0381,q0381,q0351),
       X0382(x0382,q0382,q0352),
       X0383(x0383,q0383,q0353),
       X0384(x0384,q0384,q0354),
       X0385(x0385,q0385,q0355),
       X0386(x0386,q0386,q0356),
       X0387(x0387,q0387,q0357),
       X0388(x0388,q0388,q0358),
       X0389(x0389,q0389,q0359),
       X0390(x0390,q0390,q0360);

and    A0361(a0361,n0331,o3130,q11_1,oms),
       A0362(a0362,x0332,o3130,q11_1,oms),
       A0363(a0363,x0333,o3130,q11_1,oms),
       A0364(a0364,x0334,o3130,q11_1,oms),
       A0365(a0365,x0335,o3130,q11_1,oms),
       A0366(a0366,x0336,o3130,q11_1,oms),
       A0367(a0367,x0337,o3130,q11_1,oms),
       A0368(a0368,x0338,o3130,q11_1,oms),
       A0369(a0369,x0339,o3130,q11_1,oms),
       A0370(a0370,x0340,o3130,q11_1,oms),
       A0371(a0371,x0341,o3130,q11_1,oms),
       A0372(a0372,x0342,o3130,q11_1,oms),
       A0373(a0373,x0343,o3130,q11_1,oms),
       A0374(a0374,x0344,o3130,q11_1,oms),
       A0375(a0375,x0345,o3130,q11_1,oms),
       A0376(a0376,x0346,o3130,q11_1,oms),
       A0377(a0377,x0347,o3130,q11_1,oms),
       A0378(a0378,x0348,o3130,q11_1,oms),
       A0379(a0379,x0349,o3130,q11_1,oms),
       A0380(a0380,x0350,o3130,q11_1,oms),
       A0381(a0381,x0351,o3130,q11_1,oms),
       A0382(a0382,x0352,o3130,q11_1,oms),
       A0383(a0383,x0353,o3130,q11_1,oms),
       A0384(a0384,x0354,o3130,q11_1,oms),
       A0385(a0385,x0355,o3130,q11_1,oms),
       A0386(a0386,x0356,o3130,q11_1,oms),
       A0387(a0387,x0357,o3130,q11_1,oms),
       A0388(a0388,x0358,o3130,q11_1,oms),
       A0389(a0389,x0359,o3130,q11_1,oms),
       A0390(a0390,x0360,o3130,q11_1,oms);

or     H036101(h036101,h036111,h036112,n1),
       H036201(h036201,h036211,h036212,n1),
       H036301(h036301,h036311,h036312,n1),
       H036401(h036401,h036411,h036412,n1),
       H036501(h036501,h036511,h036512,n1),
       H036601(h036601,h036611,h036612,n1),
       H036701(h036701,h036711,h036712,n1),
       H036801(h036801,h036811,h036812,n1),
       H036901(h036901,h036911,h036912,n1),
       H037001(h037001,h037011,h037012,n1),
       H037101(h037101,h037111,h037112,n1),
       H037201(h037201,h037211,h037212,n1),
       H037301(h037301,h037311,h037312,n1),
       H037401(h037401,h037411,h037412,n1),
       H037501(h037501,h037511,h037512,n1),
       H037601(h037601,h037611,h037612,n1),
       H037701(h037701,h037711,h037712,n1),
       H037801(h037801,h037811,h037812,n1),
       H037901(h037901,h037911,h037912,n1),
       H038001(h038001,h038011,h038012,n1),
       H038101(h038101,h038111,h038112,n1),
       H038201(h038201,h038211,h038212,n1),
       H038301(h038301,h038311,h038312,n1),
       H038401(h038401,h038411,h038412,n1),
       H038501(h038501,h038511,h038512,n1),
       H038601(h038601,h038611,h038612,n1),
       H038701(h038701,h038711,h038712,n1),
       H038801(h038801,h038811,h038812,n1),
       H038901(h038901,h038911,h038912,n1),
       H039001(h039001,h039011,h039012,n1);

and    H036111(h036111,oms0,dbv1),
       H036112(h036112,oms1,dbv1),
       H036211(h036211,oms0,dbv1),
       H036212(h036212,oms1,dbv1),
       H036311(h036311,oms0,dbv1),
       H036312(h036312,oms1,dbv1),
       H036411(h036411,oms0,dbv1),
       H036412(h036412,oms1,dbv1),
       H036511(h036511,oms0,dbv1),
       H036512(h036512,oms1,dbv1),
       H036611(h036611,oms0,dbv1),
       H036612(h036612,oms1,dbv1),
       H036711(h036711,oms0,dbv1),
       H036712(h036712,oms1,dbv1),
       H036811(h036811,oms0,dbv1),
       H036812(h036812,oms1,dbv1),
       H036911(h036911,oms0,dbv0),
       H036912(h036912,oms1,dbv0),
       H037011(h037011,oms0,dbv1),
       H037012(h037012,oms1,dbv0),
       H037111(h037111,oms0,dbv0),
       H037112(h037112,oms1,dbv1),
       H037211(h037211,oms0,dbv1),
       H037212(h037212,oms1,dbv0),
       H037311(h037311,oms0,dbv0),
       H037312(h037312,oms1,dbv1),
       H037411(h037411,oms0,dbv1),
       H037412(h037412,oms1,dbv0),
       H037511(h037511,oms0,dbv0),
       H037512(h037512,oms1,dbv0),
       H037611(h037611,oms0,dbv0),
       H037612(h037612,oms1,dbv1),
       H037711(h037711,oms0,dbv1),
       H037712(h037712,oms1,dbv0),
       H037811(h037811,oms0,dbv0),
       H037812(h037812,oms1,dbv0),
       H037911(h037911,oms0,dbv0),
       H037912(h037912,oms1,dbv0),
       H038011(h038011,oms0,dbv0),
       H038012(h038012,oms1,dbv0),
       H038111(h038111,oms0,dbv0),
       H038112(h038112,oms1,dbv0),
       H038211(h038211,oms0,dbv0),
       H038212(h038212,oms1,dbv0),
       H038311(h038311,oms0,dbv0),
       H038312(h038312,oms1,dbv0),
       H038411(h038411,oms0,dbv0),
       H038412(h038412,oms1,dbv0),
       H038511(h038511,oms0,dbv0),
       H038512(h038512,oms1,dbv0),
       H038611(h038611,oms0,dbv0),
       H038612(h038612,oms1,dbv0),
       H038711(h038711,oms0,dbv0),
       H038712(h038712,oms1,dbv0),
       H038811(h038811,oms0,dbv0),
       H038812(h038812,oms1,dbv0),
       H038911(h038911,oms0,dbv0),
       H038912(h038912,oms1,dbv0),
       H039011(h039011,oms0,dbv0),
       H039012(h039012,oms1,dbv0);
/*
not    H030121(h030121,h030102),
       H030221(h030221,h030202),
       H030321(h030321,h030302),
       H030421(h030421,h030402),
       H030521(h030521,h030502),
       H030621(h030621,h030602),
       H030721(h030721,h030702),
       H030821(h030821,h030802),
       H030921(h030921,h030902),
       H031021(h031021,h031002),
       H031121(h031121,h031102),
       H031221(h031221,h031202),
       H031321(h031321,h031302),
       H031421(h031421,h031402),
       H031521(h031521,h031502),
       H031621(h031621,h031602),
       H031721(h031721,h031702),
       H031821(h031821,h031802),
       H031921(h031921,h031902),
       H032021(h032021,h032002),
       H032121(h032121,h032102),
       H032221(h032221,h032202),
       H032321(h032321,h032302),
       H032421(h032421,h032402),
       H032521(h032521,h032502),
       H032621(h032621,h032602),
       H032721(h032721,h032702),
       H032821(h032821,h032802),
       H032921(h032921,h032902),
       H033021(h033021,h033002);
*/
or     O3130(o3130,x0361,x0362,x0363,x0364,x0365,x0366,x0367,x0368,x0369,x0370,x0371,x0372,x0373,x0374,x0375,x0376,x0377,x0378,x0379,x0380,x0381,x0382,x0383,x0384,x0385,x0386,x0387,x0388,x0389,x0390);
not    N3130(n3130,o3130);

or     H100_0(h100_0,h100_011,h100_012),
       H101_0(h101_0,h101_011,h101_012),
       H162_0(h162_0,h162_011,h162_012),
       H163_0(h163_0,h163_011,h163_012),
       H100_1(h100_1,h100_111,h100_112),
       H101_1(h101_1,h101_111,h101_112),
       H162_1(h162_1,h162_111,h162_112),
       H163_1(h163_1,h163_111,h163_112),
       H200_0(h200_0,h200_011,h200_012),
       H201_0(h201_0,h201_011,h201_012),
       H262_0(h262_0,h262_011,h262_012),
       H263_0(h263_0,h263_011,h263_012),
       H200_1(h200_1,h200_111,h200_112),
       H201_1(h201_1,h201_111,h201_112),
       H262_1(h262_1,h262_111,h262_112),
       H263_1(h263_1,h263_111,h263_112);

and    H100_011(h100_011,n1111111_1,q100_0,s1),
       H101_011(h101_011,n1111111_1,q101_0,s1),
       H162_011(h162_011,n1111111_1,q162_0,s1),
       H163_011(h163_011,n1111111_1,q163_0,s1),
       H100_012(h100_012,q1111111_1,n100_1,s1),
       H101_012(h101_012,q1111111_1,x101_1,s1),
       H162_012(h162_012,q1111111_1,x162_1,s1),
       H163_012(h163_012,q1111111_1,x163_1,s1),
       H100_111(h100_111,n1111111_1,q100_0,s1),
       H101_111(h101_111,n1111111_1,q101_0,s1),
       H162_111(h162_111,n1111111_1,q162_0,s1),
       H163_111(h163_111,n1111111_1,q163_0,s1),
       H100_112(h100_112,q1111111_1,q100_1,s1),
       H101_112(h101_112,q1111111_1,q101_1,s1),
       H162_112(h162_112,q1111111_1,q162_1,s1),
       H163_112(h163_112,q1111111_1,q163_1,s1),
       H200_011(h200_011,n0000000_1,q200_0,s1),
       H201_011(h201_011,n0000000_1,q201_0,s1),
       H262_011(h262_011,n0000000_1,q262_0,s1),
       H263_011(h263_011,n0000000_1,q263_0,s1),
       H200_012(h200_012,q0000000_1,n200_1,s1),
       H201_012(h201_012,q0000000_1,x201_1,s1),
       H262_012(h262_012,q0000000_1,x262_1,s1),
       H263_012(h263_012,q0000000_1,x263_1,s1),
       H200_111(h200_111,n0000000_1,q200_0,s1),
       H201_111(h201_111,n0000000_1,q201_0,s1),
       H262_111(h262_111,n0000000_1,q262_0,s1),
       H263_111(h263_111,n0000000_1,q263_0,s1),
       H200_112(h200_112,q0000000_1,q200_1,s1),
       H201_112(h201_112,q0000000_1,q201_1,s1),
       H262_112(h262_112,q0000000_1,q262_1,s1),
       H263_112(h263_112,q0000000_1,q263_1,s1);

or     H102_0(h102_0,h102_011,h102_012,h102_013),
       H103_0(h103_0,h103_011,h103_012,h103_013),
       H104_0(h104_0,h104_011,h104_012,h104_013),
       H105_0(h105_0,h105_011,h105_012,h105_013),
       H106_0(h106_0,h106_011,h106_012,h106_013),
       H107_0(h107_0,h107_011,h107_012,h107_013),
       H108_0(h108_0,h108_011,h108_012,h108_013),
       H109_0(h109_0,h109_011,h109_012,h109_013),
       H110_0(h110_0,h110_011,h110_012,h110_013),
       H111_0(h111_0,h111_011,h111_012,h111_013),
       H112_0(h112_0,h112_011,h112_012,h112_013),
       H113_0(h113_0,h113_011,h113_012,h113_013),
       H114_0(h114_0,h114_011,h114_012,h114_013),
       H115_0(h115_0,h115_011,h115_012,h115_013),
       H116_0(h116_0,h116_011,h116_012,h116_013),
       H117_0(h117_0,h117_011,h117_012,h117_013),
       H118_0(h118_0,h118_011,h118_012,h118_013),
       H119_0(h119_0,h119_011,h119_012,h119_013),
       H120_0(h120_0,h120_011,h120_012,h120_013),
       H121_0(h121_0,h121_011,h121_012,h121_013),
       H122_0(h122_0,h122_011,h122_012,h122_013),
       H123_0(h123_0,h123_011,h123_012,h123_013),
       H124_0(h124_0,h124_011,h124_012,h124_013),
       H125_0(h125_0,h125_011,h125_012,h125_013),
       H126_0(h126_0,h126_011,h126_012,h126_013),
       H127_0(h127_0,h127_011,h127_012,h127_013),
       H128_0(h128_0,h128_011,h128_012,h128_013),
       H129_0(h129_0,h129_011,h129_012,h129_013),
       H130_0(h130_0,h130_011,h130_012,h130_013),
       H131_0(h131_0,h131_011,h131_012,h131_013),
       H132_0(h132_0,h132_011,h132_012,h132_013),
       H133_0(h133_0,h133_011,h133_012,h133_013),
       H134_0(h134_0,h134_011,h134_012,h134_013),
       H135_0(h135_0,h135_011,h135_012,h135_013),
       H136_0(h136_0,h136_011,h136_012,h136_013),
       H137_0(h137_0,h137_011,h137_012,h137_013),
       H138_0(h138_0,h138_011,h138_012,h138_013),
       H139_0(h139_0,h139_011,h139_012,h139_013),
       H140_0(h140_0,h140_011,h140_012,h140_013),
       H141_0(h141_0,h141_011,h141_012,h141_013),
       H142_0(h142_0,h142_011,h142_012,h142_013),
       H143_0(h143_0,h143_011,h143_012,h143_013),
       H144_0(h144_0,h144_011,h144_012,h144_013),
       H145_0(h145_0,h145_011,h145_012,h145_013),
       H146_0(h146_0,h146_011,h146_012,h146_013),
       H147_0(h147_0,h147_011,h147_012,h147_013),
       H148_0(h148_0,h148_011,h148_012,h148_013),
       H149_0(h149_0,h149_011,h149_012,h149_013),
       H150_0(h150_0,h150_011,h150_012,h150_013),
       H151_0(h151_0,h151_011,h151_012,h151_013),
       H152_0(h152_0,h152_011,h152_012,h152_013),
       H153_0(h153_0,h153_011,h153_012,h153_013),
       H154_0(h154_0,h154_011,h154_012,h154_013),
       H155_0(h155_0,h155_011,h155_012,h155_013),
       H156_0(h156_0,h156_011,h156_012,h156_013),
       H157_0(h157_0,h157_011,h157_012,h157_013),
       H158_0(h158_0,h158_011,h158_012,h158_013),
       H159_0(h159_0,h159_011,h159_012,h159_013),
       H160_0(h160_0,h160_011,h160_012,h160_013),
       H161_0(h161_0,h161_011,h161_012,h161_013),
       H102_1(h102_1,h102_111,h102_112),
       H103_1(h103_1,h103_111,h103_112),
       H104_1(h104_1,h104_111,h104_112),
       H105_1(h105_1,h105_111,h105_112),
       H106_1(h106_1,h106_111,h106_112),
       H107_1(h107_1,h107_111,h107_112),
       H108_1(h108_1,h108_111,h108_112),
       H109_1(h109_1,h109_111,h109_112),
       H110_1(h110_1,h110_111,h110_112),
       H111_1(h111_1,h111_111,h111_112),
       H112_1(h112_1,h112_111,h112_112),
       H113_1(h113_1,h113_111,h113_112),
       H114_1(h114_1,h114_111,h114_112),
       H115_1(h115_1,h115_111,h115_112),
       H116_1(h116_1,h116_111,h116_112),
       H117_1(h117_1,h117_111,h117_112),
       H118_1(h118_1,h118_111,h118_112),
       H119_1(h119_1,h119_111,h119_112),
       H120_1(h120_1,h120_111,h120_112),
       H121_1(h121_1,h121_111,h121_112),
       H122_1(h122_1,h122_111,h122_112),
       H123_1(h123_1,h123_111,h123_112),
       H124_1(h124_1,h124_111,h124_112),
       H125_1(h125_1,h125_111,h125_112),
       H126_1(h126_1,h126_111,h126_112),
       H127_1(h127_1,h127_111,h127_112),
       H128_1(h128_1,h128_111,h128_112),
       H129_1(h129_1,h129_111,h129_112),
       H130_1(h130_1,h130_111,h130_112),
       H131_1(h131_1,h131_111,h131_112),
       H132_1(h132_1,h132_111,h132_112),
       H133_1(h133_1,h133_111,h133_112),
       H134_1(h134_1,h134_111,h134_112),
       H135_1(h135_1,h135_111,h135_112),
       H136_1(h136_1,h136_111,h136_112),
       H137_1(h137_1,h137_111,h137_112),
       H138_1(h138_1,h138_111,h138_112),
       H139_1(h139_1,h139_111,h139_112),
       H140_1(h140_1,h140_111,h140_112),
       H141_1(h141_1,h141_111,h141_112),
       H142_1(h142_1,h142_111,h142_112),
       H143_1(h143_1,h143_111,h143_112),
       H144_1(h144_1,h144_111,h144_112),
       H145_1(h145_1,h145_111,h145_112),
       H146_1(h146_1,h146_111,h146_112),
       H147_1(h147_1,h147_111,h147_112),
       H148_1(h148_1,h148_111,h148_112),
       H149_1(h149_1,h149_111,h149_112),
       H150_1(h150_1,h150_111,h150_112),
       H151_1(h151_1,h151_111,h151_112),
       H152_1(h152_1,h152_111,h152_112),
       H153_1(h153_1,h153_111,h153_112),
       H154_1(h154_1,h154_111,h154_112),
       H155_1(h155_1,h155_111,h155_112),
       H156_1(h156_1,h156_111,h156_112),
       H157_1(h157_1,h157_111,h157_112),
       H158_1(h158_1,h158_111,h158_112),
       H159_1(h159_1,h159_111,h159_112),
       H160_1(h160_1,h160_111,h160_112),
       H161_1(h161_1,h161_111,h161_112),
       H202_0(h202_0,h202_011,h202_012,h202_013),
       H203_0(h203_0,h203_011,h203_012,h203_013),
       H204_0(h204_0,h204_011,h204_012,h204_013),
       H205_0(h205_0,h205_011,h205_012,h205_013),
       H206_0(h206_0,h206_011,h206_012,h206_013),
       H207_0(h207_0,h207_011,h207_012,h207_013),
       H208_0(h208_0,h208_011,h208_012,h208_013),
       H209_0(h209_0,h209_011,h209_012,h209_013),
       H210_0(h210_0,h210_011,h210_012,h210_013),
       H211_0(h211_0,h211_011,h211_012,h211_013),
       H212_0(h212_0,h212_011,h212_012,h212_013),
       H213_0(h213_0,h213_011,h213_012,h213_013),
       H214_0(h214_0,h214_011,h214_012,h214_013),
       H215_0(h215_0,h215_011,h215_012,h215_013),
       H216_0(h216_0,h216_011,h216_012,h216_013),
       H217_0(h217_0,h217_011,h217_012,h217_013),
       H218_0(h218_0,h218_011,h218_012,h218_013),
       H219_0(h219_0,h219_011,h219_012,h219_013),
       H220_0(h220_0,h220_011,h220_012,h220_013),
       H221_0(h221_0,h221_011,h221_012,h221_013),
       H222_0(h222_0,h222_011,h222_012,h222_013),
       H223_0(h223_0,h223_011,h223_012,h223_013),
       H224_0(h224_0,h224_011,h224_012,h224_013),
       H225_0(h225_0,h225_011,h225_012,h225_013),
       H226_0(h226_0,h226_011,h226_012,h226_013),
       H227_0(h227_0,h227_011,h227_012,h227_013),
       H228_0(h228_0,h228_011,h228_012,h228_013),
       H229_0(h229_0,h229_011,h229_012,h229_013),
       H230_0(h230_0,h230_011,h230_012,h230_013),
       H231_0(h231_0,h231_011,h231_012,h231_013),
       H232_0(h232_0,h232_011,h232_012,h232_013),
       H233_0(h233_0,h233_011,h233_012,h233_013),
       H234_0(h234_0,h234_011,h234_012,h234_013),
       H235_0(h235_0,h235_011,h235_012,h235_013),
       H236_0(h236_0,h236_011,h236_012,h236_013),
       H237_0(h237_0,h237_011,h237_012,h237_013),
       H238_0(h238_0,h238_011,h238_012,h238_013),
       H239_0(h239_0,h239_011,h239_012,h239_013),
       H240_0(h240_0,h240_011,h240_012,h240_013),
       H241_0(h241_0,h241_011,h241_012,h241_013),
       H242_0(h242_0,h242_011,h242_012,h242_013),
       H243_0(h243_0,h243_011,h243_012,h243_013),
       H244_0(h244_0,h244_011,h244_012,h244_013),
       H245_0(h245_0,h245_011,h245_012,h245_013),
       H246_0(h246_0,h246_011,h246_012,h246_013),
       H247_0(h247_0,h247_011,h247_012,h247_013),
       H248_0(h248_0,h248_011,h248_012,h248_013),
       H249_0(h249_0,h249_011,h249_012,h249_013),
       H250_0(h250_0,h250_011,h250_012,h250_013),
       H251_0(h251_0,h251_011,h251_012,h251_013),
       H252_0(h252_0,h252_011,h252_012,h252_013),
       H253_0(h253_0,h253_011,h253_012,h253_013),
       H254_0(h254_0,h254_011,h254_012,h254_013),
       H255_0(h255_0,h255_011,h255_012,h255_013),
       H256_0(h256_0,h256_011,h256_012,h256_013),
       H257_0(h257_0,h257_011,h257_012,h257_013),
       H258_0(h258_0,h258_011,h258_012,h258_013),
       H259_0(h259_0,h259_011,h259_012,h259_013),
       H260_0(h260_0,h260_011,h260_012,h260_013),
       H261_0(h261_0,h261_011,h261_012,h261_013),
       H202_1(h202_1,h202_111,h202_112),
       H203_1(h203_1,h203_111,h203_112),
       H204_1(h204_1,h204_111,h204_112),
       H205_1(h205_1,h205_111,h205_112),
       H206_1(h206_1,h206_111,h206_112),
       H207_1(h207_1,h207_111,h207_112),
       H208_1(h208_1,h208_111,h208_112),
       H209_1(h209_1,h209_111,h209_112),
       H210_1(h210_1,h210_111,h210_112),
       H211_1(h211_1,h211_111,h211_112),
       H212_1(h212_1,h212_111,h212_112),
       H213_1(h213_1,h213_111,h213_112),
       H214_1(h214_1,h214_111,h214_112),
       H215_1(h215_1,h215_111,h215_112),
       H216_1(h216_1,h216_111,h216_112),
       H217_1(h217_1,h217_111,h217_112),
       H218_1(h218_1,h218_111,h218_112),
       H219_1(h219_1,h219_111,h219_112),
       H220_1(h220_1,h220_111,h220_112),
       H221_1(h221_1,h221_111,h221_112),
       H222_1(h222_1,h222_111,h222_112),
       H223_1(h223_1,h223_111,h223_112),
       H224_1(h224_1,h224_111,h224_112),
       H225_1(h225_1,h225_111,h225_112),
       H226_1(h226_1,h226_111,h226_112),
       H227_1(h227_1,h227_111,h227_112),
       H228_1(h228_1,h228_111,h228_112),
       H229_1(h229_1,h229_111,h229_112),
       H230_1(h230_1,h230_111,h230_112),
       H231_1(h231_1,h231_111,h231_112),
       H232_1(h232_1,h232_111,h232_112),
       H233_1(h233_1,h233_111,h233_112),
       H234_1(h234_1,h234_111,h234_112),
       H235_1(h235_1,h235_111,h235_112),
       H236_1(h236_1,h236_111,h236_112),
       H237_1(h237_1,h237_111,h237_112),
       H238_1(h238_1,h238_111,h238_112),
       H239_1(h239_1,h239_111,h239_112),
       H240_1(h240_1,h240_111,h240_112),
       H241_1(h241_1,h241_111,h241_112),
       H242_1(h242_1,h242_111,h242_112),
       H243_1(h243_1,h243_111,h243_112),
       H244_1(h244_1,h244_111,h244_112),
       H245_1(h245_1,h245_111,h245_112),
       H246_1(h246_1,h246_111,h246_112),
       H247_1(h247_1,h247_111,h247_112),
       H248_1(h248_1,h248_111,h248_112),
       H249_1(h249_1,h249_111,h249_112),
       H250_1(h250_1,h250_111,h250_112),
       H251_1(h251_1,h251_111,h251_112),
       H252_1(h252_1,h252_111,h252_112),
       H253_1(h253_1,h253_111,h253_112),
       H254_1(h254_1,h254_111,h254_112),
       H255_1(h255_1,h255_111,h255_112),
       H256_1(h256_1,h256_111,h256_112),
       H257_1(h257_1,h257_111,h257_112),
       H258_1(h258_1,h258_111,h258_112),
       H259_1(h259_1,h259_111,h259_112),
       H260_1(h260_1,h260_111,h260_112),
       H261_1(h261_1,h261_111,h261_112);

and    H102_011(h102_011,o5110,q102_0),
       H103_011(h103_011,o5110,q103_0),
       H104_011(h104_011,o5110,q104_0),
       H105_011(h105_011,o5110,q105_0),
       H106_011(h106_011,o5110,q106_0),
       H107_011(h107_011,o5110,q107_0),
       H108_011(h108_011,o5110,q108_0),
       H109_011(h109_011,o5110,q109_0),
       H110_011(h110_011,o5110,q110_0),
       H111_011(h111_011,o5110,q111_0),
       H112_011(h112_011,o5110,q112_0),
       H113_011(h113_011,o5110,q113_0),
       H114_011(h114_011,o5110,q114_0),
       H115_011(h115_011,o5110,q115_0),
       H116_011(h116_011,o5110,q116_0),
       H117_011(h117_011,o5110,q117_0),
       H118_011(h118_011,o5110,q118_0),
       H119_011(h119_011,o5110,q119_0),
       H120_011(h120_011,o5110,q120_0),
       H121_011(h121_011,o5110,q121_0),
       H122_011(h122_011,o5110,q122_0),
       H123_011(h123_011,o5110,q123_0),
       H124_011(h124_011,o5110,q124_0),
       H125_011(h125_011,o5110,q125_0),
       H126_011(h126_011,o5110,q126_0),
       H127_011(h127_011,o5110,q127_0),
       H128_011(h128_011,o5110,q128_0),
       H129_011(h129_011,o5110,q129_0),
       H130_011(h130_011,o5110,q130_0),
       H131_011(h131_011,o5110,q131_0),
       H132_011(h132_011,o5110,q132_0),
       H133_011(h133_011,o5110,q133_0),
       H134_011(h134_011,o5110,q134_0),
       H135_011(h135_011,o5110,q135_0),
       H136_011(h136_011,o5110,q136_0),
       H137_011(h137_011,o5110,q137_0),
       H138_011(h138_011,o5110,q138_0),
       H139_011(h139_011,o5110,q139_0),
       H140_011(h140_011,o5110,q140_0),
       H141_011(h141_011,o5110,q141_0),
       H142_011(h142_011,o5110,q142_0),
       H143_011(h143_011,o5110,q143_0),
       H144_011(h144_011,o5110,q144_0),
       H145_011(h145_011,o5110,q145_0),
       H146_011(h146_011,o5110,q146_0),
       H147_011(h147_011,o5110,q147_0),
       H148_011(h148_011,o5110,q148_0),
       H149_011(h149_011,o5110,q149_0),
       H150_011(h150_011,o5110,q150_0),
       H151_011(h151_011,o5110,q151_0),
       H152_011(h152_011,o5110,q152_0),
       H153_011(h153_011,o5110,q153_0),
       H154_011(h154_011,o5110,q154_0),
       H155_011(h155_011,o5110,q155_0),
       H156_011(h156_011,o5110,q156_0),
       H157_011(h157_011,o5110,q157_0),
       H158_011(h158_011,o5110,q158_0),
       H159_011(h159_011,o5110,q159_0),
       H160_011(h160_011,o5110,q160_0),
       H161_011(h161_011,o5110,q161_0),
       H102_012(h102_012,n5110,sl,q161_1),
       H103_012(h103_012,n5110,sl,q102_1),
       H104_012(h104_012,n5110,sl,q103_1),
       H105_012(h105_012,n5110,sl,q104_1),
       H106_012(h106_012,n5110,sl,q105_1),
       H107_012(h107_012,n5110,sl,q106_1),
       H108_012(h108_012,n5110,sl,q107_1),
       H109_012(h109_012,n5110,sl,q108_1),
       H110_012(h110_012,n5110,sl,q109_1),
       H111_012(h111_012,n5110,sl,q110_1),
       H112_012(h112_012,n5110,sl,q111_1),
       H113_012(h113_012,n5110,sl,q112_1),
       H114_012(h114_012,n5110,sl,q113_1),
       H115_012(h115_012,n5110,sl,q114_1),
       H116_012(h116_012,n5110,sl,q115_1),
       H117_012(h117_012,n5110,sl,q116_1),
       H118_012(h118_012,n5110,sl,q117_1),
       H119_012(h119_012,n5110,sl,q118_1),
       H120_012(h120_012,n5110,sl,q119_1),
       H121_012(h121_012,n5110,sl,q120_1),
       H122_012(h122_012,n5110,sl,q121_1),
       H123_012(h123_012,n5110,sl,q122_1),
       H124_012(h124_012,n5110,sl,q123_1),
       H125_012(h125_012,n5110,sl,q124_1),
       H126_012(h126_012,n5110,sl,q125_1),
       H127_012(h127_012,n5110,sl,q126_1),
       H128_012(h128_012,n5110,sl,q127_1),
       H129_012(h129_012,n5110,sl,q128_1),
       H130_012(h130_012,n5110,sl,q129_1),
       H131_012(h131_012,n5110,sl,q130_1),
       H132_012(h132_012,n5110,sl,q131_1),
       H133_012(h133_012,n5110,sl,q132_1),
       H134_012(h134_012,n5110,sl,q133_1),
       H135_012(h135_012,n5110,sl,q134_1),
       H136_012(h136_012,n5110,sl,q135_1),
       H137_012(h137_012,n5110,sl,q136_1),
       H138_012(h138_012,n5110,sl,q137_1),
       H139_012(h139_012,n5110,sl,q138_1),
       H140_012(h140_012,n5110,sl,q139_1),
       H141_012(h141_012,n5110,sl,q140_1),
       H142_012(h142_012,n5110,sl,q141_1),
       H143_012(h143_012,n5110,sl,q142_1),
       H144_012(h144_012,n5110,sl,q143_1),
       H145_012(h145_012,n5110,sl,q144_1),
       H146_012(h146_012,n5110,sl,q145_1),
       H147_012(h147_012,n5110,sl,q146_1),
       H148_012(h148_012,n5110,sl,q147_1),
       H149_012(h149_012,n5110,sl,q148_1),
       H150_012(h150_012,n5110,sl,q149_1),
       H151_012(h151_012,n5110,sl,q150_1),
       H152_012(h152_012,n5110,sl,q151_1),
       H153_012(h153_012,n5110,sl,q152_1),
       H154_012(h154_012,n5110,sl,q153_1),
       H155_012(h155_012,n5110,sl,q154_1),
       H156_012(h156_012,n5110,sl,q155_1),
       H157_012(h157_012,n5110,sl,q156_1),
       H158_012(h158_012,n5110,sl,q157_1),
       H159_012(h159_012,n5110,sl,q158_1),
       H160_012(h160_012,n5110,sl,q159_1),
       H161_012(h161_012,n5110,sl,q160_1),
       H102_013(h102_013,n5110,sr,q103_1),
       H103_013(h103_013,n5110,sr,q104_1),
       H104_013(h104_013,n5110,sr,q105_1),
       H105_013(h105_013,n5110,sr,q106_1),
       H106_013(h106_013,n5110,sr,q107_1),
       H107_013(h107_013,n5110,sr,q108_1),
       H108_013(h108_013,n5110,sr,q109_1),
       H109_013(h109_013,n5110,sr,q110_1),
       H110_013(h110_013,n5110,sr,q111_1),
       H111_013(h111_013,n5110,sr,q112_1),
       H112_013(h112_013,n5110,sr,q113_1),
       H113_013(h113_013,n5110,sr,q114_1),
       H114_013(h114_013,n5110,sr,q115_1),
       H115_013(h115_013,n5110,sr,q116_1),
       H116_013(h116_013,n5110,sr,q117_1),
       H117_013(h117_013,n5110,sr,q118_1),
       H118_013(h118_013,n5110,sr,q119_1),
       H119_013(h119_013,n5110,sr,q120_1),
       H120_013(h120_013,n5110,sr,q121_1),
       H121_013(h121_013,n5110,sr,q122_1),
       H122_013(h122_013,n5110,sr,q123_1),
       H123_013(h123_013,n5110,sr,q124_1),
       H124_013(h124_013,n5110,sr,q125_1),
       H125_013(h125_013,n5110,sr,q126_1),
       H126_013(h126_013,n5110,sr,q127_1),
       H127_013(h127_013,n5110,sr,q128_1),
       H128_013(h128_013,n5110,sr,q129_1),
       H129_013(h129_013,n5110,sr,q130_1),
       H130_013(h130_013,n5110,sr,q131_1),
       H131_013(h131_013,n5110,sr,q132_1),
       H132_013(h132_013,n5110,sr,q133_1),
       H133_013(h133_013,n5110,sr,q134_1),
       H134_013(h134_013,n5110,sr,q135_1),
       H135_013(h135_013,n5110,sr,q136_1),
       H136_013(h136_013,n5110,sr,q137_1),
       H137_013(h137_013,n5110,sr,q138_1),
       H138_013(h138_013,n5110,sr,q139_1),
       H139_013(h139_013,n5110,sr,q140_1),
       H140_013(h140_013,n5110,sr,q141_1),
       H141_013(h141_013,n5110,sr,q142_1),
       H142_013(h142_013,n5110,sr,q143_1),
       H143_013(h143_013,n5110,sr,q144_1),
       H144_013(h144_013,n5110,sr,q145_1),
       H145_013(h145_013,n5110,sr,q146_1),
       H146_013(h146_013,n5110,sr,q147_1),
       H147_013(h147_013,n5110,sr,q148_1),
       H148_013(h148_013,n5110,sr,q149_1),
       H149_013(h149_013,n5110,sr,q150_1),
       H150_013(h150_013,n5110,sr,q151_1),
       H151_013(h151_013,n5110,sr,q152_1),
       H152_013(h152_013,n5110,sr,q153_1),
       H153_013(h153_013,n5110,sr,q154_1),
       H154_013(h154_013,n5110,sr,q155_1),
       H155_013(h155_013,n5110,sr,q156_1),
       H156_013(h156_013,n5110,sr,q157_1),
       H157_013(h157_013,n5110,sr,q158_1),
       H158_013(h158_013,n5110,sr,q159_1),
       H159_013(h159_013,n5110,sr,q160_1),
       H160_013(h160_013,n5110,sr,q161_1),
       H161_013(h161_013,n5110,sr,q102_1),
       H102_111(h102_111,o5110,q102_0),
       H103_111(h103_111,o5110,q103_0),
       H104_111(h104_111,o5110,q104_0),
       H105_111(h105_111,o5110,q105_0),
       H106_111(h106_111,o5110,q106_0),
       H107_111(h107_111,o5110,q107_0),
       H108_111(h108_111,o5110,q108_0),
       H109_111(h109_111,o5110,q109_0),
       H110_111(h110_111,o5110,q110_0),
       H111_111(h111_111,o5110,q111_0),
       H112_111(h112_111,o5110,q112_0),
       H113_111(h113_111,o5110,q113_0),
       H114_111(h114_111,o5110,q114_0),
       H115_111(h115_111,o5110,q115_0),
       H116_111(h116_111,o5110,q116_0),
       H117_111(h117_111,o5110,q117_0),
       H118_111(h118_111,o5110,q118_0),
       H119_111(h119_111,o5110,q119_0),
       H120_111(h120_111,o5110,q120_0),
       H121_111(h121_111,o5110,q121_0),
       H122_111(h122_111,o5110,q122_0),
       H123_111(h123_111,o5110,q123_0),
       H124_111(h124_111,o5110,q124_0),
       H125_111(h125_111,o5110,q125_0),
       H126_111(h126_111,o5110,q126_0),
       H127_111(h127_111,o5110,q127_0),
       H128_111(h128_111,o5110,q128_0),
       H129_111(h129_111,o5110,q129_0),
       H130_111(h130_111,o5110,q130_0),
       H131_111(h131_111,o5110,q131_0),
       H132_111(h132_111,o5110,q132_0),
       H133_111(h133_111,o5110,q133_0),
       H134_111(h134_111,o5110,q134_0),
       H135_111(h135_111,o5110,q135_0),
       H136_111(h136_111,o5110,q136_0),
       H137_111(h137_111,o5110,q137_0),
       H138_111(h138_111,o5110,q138_0),
       H139_111(h139_111,o5110,q139_0),
       H140_111(h140_111,o5110,q140_0),
       H141_111(h141_111,o5110,q141_0),
       H142_111(h142_111,o5110,q142_0),
       H143_111(h143_111,o5110,q143_0),
       H144_111(h144_111,o5110,q144_0),
       H145_111(h145_111,o5110,q145_0),
       H146_111(h146_111,o5110,q146_0),
       H147_111(h147_111,o5110,q147_0),
       H148_111(h148_111,o5110,q148_0),
       H149_111(h149_111,o5110,q149_0),
       H150_111(h150_111,o5110,q150_0),
       H151_111(h151_111,o5110,q151_0),
       H152_111(h152_111,o5110,q152_0),
       H153_111(h153_111,o5110,q153_0),
       H154_111(h154_111,o5110,q154_0),
       H155_111(h155_111,o5110,q155_0),
       H156_111(h156_111,o5110,q156_0),
       H157_111(h157_111,o5110,q157_0),
       H158_111(h158_111,o5110,q158_0),
       H159_111(h159_111,o5110,q159_0),
       H160_111(h160_111,o5110,q160_0),
       H161_111(h161_111,o5110,q161_0),
       H102_112(h102_112,n5110,q102_1),
       H103_112(h103_112,n5110,q103_1),
       H104_112(h104_112,n5110,q104_1),
       H105_112(h105_112,n5110,q105_1),
       H106_112(h106_112,n5110,q106_1),
       H107_112(h107_112,n5110,q107_1),
       H108_112(h108_112,n5110,q108_1),
       H109_112(h109_112,n5110,q109_1),
       H110_112(h110_112,n5110,q110_1),
       H111_112(h111_112,n5110,q111_1),
       H112_112(h112_112,n5110,q112_1),
       H113_112(h113_112,n5110,q113_1),
       H114_112(h114_112,n5110,q114_1),
       H115_112(h115_112,n5110,q115_1),
       H116_112(h116_112,n5110,q116_1),
       H117_112(h117_112,n5110,q117_1),
       H118_112(h118_112,n5110,q118_1),
       H119_112(h119_112,n5110,q119_1),
       H120_112(h120_112,n5110,q120_1),
       H121_112(h121_112,n5110,q121_1),
       H122_112(h122_112,n5110,q122_1),
       H123_112(h123_112,n5110,q123_1),
       H124_112(h124_112,n5110,q124_1),
       H125_112(h125_112,n5110,q125_1),
       H126_112(h126_112,n5110,q126_1),
       H127_112(h127_112,n5110,q127_1),
       H128_112(h128_112,n5110,q128_1),
       H129_112(h129_112,n5110,q129_1),
       H130_112(h130_112,n5110,q130_1),
       H131_112(h131_112,n5110,q131_1),
       H132_112(h132_112,n5110,q132_1),
       H133_112(h133_112,n5110,q133_1),
       H134_112(h134_112,n5110,q134_1),
       H135_112(h135_112,n5110,q135_1),
       H136_112(h136_112,n5110,q136_1),
       H137_112(h137_112,n5110,q137_1),
       H138_112(h138_112,n5110,q138_1),
       H139_112(h139_112,n5110,q139_1),
       H140_112(h140_112,n5110,q140_1),
       H141_112(h141_112,n5110,q141_1),
       H142_112(h142_112,n5110,q142_1),
       H143_112(h143_112,n5110,q143_1),
       H144_112(h144_112,n5110,q144_1),
       H145_112(h145_112,n5110,q145_1),
       H146_112(h146_112,n5110,q146_1),
       H147_112(h147_112,n5110,q147_1),
       H148_112(h148_112,n5110,q148_1),
       H149_112(h149_112,n5110,q149_1),
       H150_112(h150_112,n5110,q150_1),
       H151_112(h151_112,n5110,q151_1),
       H152_112(h152_112,n5110,q152_1),
       H153_112(h153_112,n5110,q153_1),
       H154_112(h154_112,n5110,q154_1),
       H155_112(h155_112,n5110,q155_1),
       H156_112(h156_112,n5110,q156_1),
       H157_112(h157_112,n5110,q157_1),
       H158_112(h158_112,n5110,q158_1),
       H159_112(h159_112,n5110,q159_1),
       H160_112(h160_112,n5110,q160_1),
       H161_112(h161_112,n5110,q161_1),
       H202_011(h202_011,o1170,q202_0),
       H203_011(h203_011,o1170,q203_0),
       H204_011(h204_011,o1170,q204_0),
       H205_011(h205_011,o1170,q205_0),
       H206_011(h206_011,o1170,q206_0),
       H207_011(h207_011,o1170,q207_0),
       H208_011(h208_011,o1170,q208_0),
       H209_011(h209_011,o1170,q209_0),
       H210_011(h210_011,o1170,q210_0),
       H211_011(h211_011,o1170,q211_0),
       H212_011(h212_011,o1170,q212_0),
       H213_011(h213_011,o1170,q213_0),
       H214_011(h214_011,o1170,q214_0),
       H215_011(h215_011,o1170,q215_0),
       H216_011(h216_011,o1170,q216_0),
       H217_011(h217_011,o1170,q217_0),
       H218_011(h218_011,o1170,q218_0),
       H219_011(h219_011,o1170,q219_0),
       H220_011(h220_011,o1170,q220_0),
       H221_011(h221_011,o1170,q221_0),
       H222_011(h222_011,o1170,q222_0),
       H223_011(h223_011,o1170,q223_0),
       H224_011(h224_011,o1170,q224_0),
       H225_011(h225_011,o1170,q225_0),
       H226_011(h226_011,o1170,q226_0),
       H227_011(h227_011,o1170,q227_0),
       H228_011(h228_011,o1170,q228_0),
       H229_011(h229_011,o1170,q229_0),
       H230_011(h230_011,o1170,q230_0),
       H231_011(h231_011,o1170,q231_0),
       H232_011(h232_011,o1170,q232_0),
       H233_011(h233_011,o1170,q233_0),
       H234_011(h234_011,o1170,q234_0),
       H235_011(h235_011,o1170,q235_0),
       H236_011(h236_011,o1170,q236_0),
       H237_011(h237_011,o1170,q237_0),
       H238_011(h238_011,o1170,q238_0),
       H239_011(h239_011,o1170,q239_0),
       H240_011(h240_011,o1170,q240_0),
       H241_011(h241_011,o1170,q241_0),
       H242_011(h242_011,o1170,q242_0),
       H243_011(h243_011,o1170,q243_0),
       H244_011(h244_011,o1170,q244_0),
       H245_011(h245_011,o1170,q245_0),
       H246_011(h246_011,o1170,q246_0),
       H247_011(h247_011,o1170,q247_0),
       H248_011(h248_011,o1170,q248_0),
       H249_011(h249_011,o1170,q249_0),
       H250_011(h250_011,o1170,q250_0),
       H251_011(h251_011,o1170,q251_0),
       H252_011(h252_011,o1170,q252_0),
       H253_011(h253_011,o1170,q253_0),
       H254_011(h254_011,o1170,q254_0),
       H255_011(h255_011,o1170,q255_0),
       H256_011(h256_011,o1170,q256_0),
       H257_011(h257_011,o1170,q257_0),
       H258_011(h258_011,o1170,q258_0),
       H259_011(h259_011,o1170,q259_0),
       H260_011(h260_011,o1170,q260_0),
       H261_011(h261_011,o1170,q261_0),
       H202_012(h202_012,n1170,kr,q261_1),
       H203_012(h203_012,n1170,kr,q202_1),
       H204_012(h204_012,n1170,kr,q203_1),
       H205_012(h205_012,n1170,kr,q204_1),
       H206_012(h206_012,n1170,kr,q205_1),
       H207_012(h207_012,n1170,kr,q206_1),
       H208_012(h208_012,n1170,kr,q207_1),
       H209_012(h209_012,n1170,kr,q208_1),
       H210_012(h210_012,n1170,kr,q209_1),
       H211_012(h211_012,n1170,kr,q210_1),
       H212_012(h212_012,n1170,kr,q211_1),
       H213_012(h213_012,n1170,kr,q212_1),
       H214_012(h214_012,n1170,kr,q213_1),
       H215_012(h215_012,n1170,kr,q214_1),
       H216_012(h216_012,n1170,kr,q215_1),
       H217_012(h217_012,n1170,kr,q216_1),
       H218_012(h218_012,n1170,kr,q217_1),
       H219_012(h219_012,n1170,kr,q218_1),
       H220_012(h220_012,n1170,kr,q219_1),
       H221_012(h221_012,n1170,kr,q220_1),
       H222_012(h222_012,n1170,kr,q221_1),
       H223_012(h223_012,n1170,kr,q222_1),
       H224_012(h224_012,n1170,kr,q223_1),
       H225_012(h225_012,n1170,kr,q224_1),
       H226_012(h226_012,n1170,kr,q225_1),
       H227_012(h227_012,n1170,kr,q226_1),
       H228_012(h228_012,n1170,kr,q227_1),
       H229_012(h229_012,n1170,kr,q228_1),
       H230_012(h230_012,n1170,kr,q229_1),
       H231_012(h231_012,n1170,kr,q230_1),
       H232_012(h232_012,n1170,kr,q231_1),
       H233_012(h233_012,n1170,kr,q232_1),
       H234_012(h234_012,n1170,kr,q233_1),
       H235_012(h235_012,n1170,kr,q234_1),
       H236_012(h236_012,n1170,kr,q235_1),
       H237_012(h237_012,n1170,kr,q236_1),
       H238_012(h238_012,n1170,kr,q237_1),
       H239_012(h239_012,n1170,kr,q238_1),
       H240_012(h240_012,n1170,kr,q239_1),
       H241_012(h241_012,n1170,kr,q240_1),
       H242_012(h242_012,n1170,kr,q241_1),
       H243_012(h243_012,n1170,kr,q242_1),
       H244_012(h244_012,n1170,kr,q243_1),
       H245_012(h245_012,n1170,kr,q244_1),
       H246_012(h246_012,n1170,kr,q245_1),
       H247_012(h247_012,n1170,kr,q246_1),
       H248_012(h248_012,n1170,kr,q247_1),
       H249_012(h249_012,n1170,kr,q248_1),
       H250_012(h250_012,n1170,kr,q249_1),
       H251_012(h251_012,n1170,kr,q250_1),
       H252_012(h252_012,n1170,kr,q251_1),
       H253_012(h253_012,n1170,kr,q252_1),
       H254_012(h254_012,n1170,kr,q253_1),
       H255_012(h255_012,n1170,kr,q254_1),
       H256_012(h256_012,n1170,kr,q255_1),
       H257_012(h257_012,n1170,kr,q256_1),
       H258_012(h258_012,n1170,kr,q257_1),
       H259_012(h259_012,n1170,kr,q258_1),
       H260_012(h260_012,n1170,kr,q259_1),
       H261_012(h261_012,n1170,kr,q260_1),
       H202_013(h202_013,n1170,kl,q203_1),
       H203_013(h203_013,n1170,kl,q204_1),
       H204_013(h204_013,n1170,kl,q205_1),
       H205_013(h205_013,n1170,kl,q206_1),
       H206_013(h206_013,n1170,kl,q207_1),
       H207_013(h207_013,n1170,kl,q208_1),
       H208_013(h208_013,n1170,kl,q209_1),
       H209_013(h209_013,n1170,kl,q210_1),
       H210_013(h210_013,n1170,kl,q211_1),
       H211_013(h211_013,n1170,kl,q212_1),
       H212_013(h212_013,n1170,kl,q213_1),
       H213_013(h213_013,n1170,kl,q214_1),
       H214_013(h214_013,n1170,kl,q215_1),
       H215_013(h215_013,n1170,kl,q216_1),
       H216_013(h216_013,n1170,kl,q217_1),
       H217_013(h217_013,n1170,kl,q218_1),
       H218_013(h218_013,n1170,kl,q219_1),
       H219_013(h219_013,n1170,kl,q220_1),
       H220_013(h220_013,n1170,kl,q221_1),
       H221_013(h221_013,n1170,kl,q222_1),
       H222_013(h222_013,n1170,kl,q223_1),
       H223_013(h223_013,n1170,kl,q224_1),
       H224_013(h224_013,n1170,kl,q225_1),
       H225_013(h225_013,n1170,kl,q226_1),
       H226_013(h226_013,n1170,kl,q227_1),
       H227_013(h227_013,n1170,kl,q228_1),
       H228_013(h228_013,n1170,kl,q229_1),
       H229_013(h229_013,n1170,kl,q230_1),
       H230_013(h230_013,n1170,kl,q231_1),
       H231_013(h231_013,n1170,kl,q232_1),
       H232_013(h232_013,n1170,kl,q233_1),
       H233_013(h233_013,n1170,kl,q234_1),
       H234_013(h234_013,n1170,kl,q235_1),
       H235_013(h235_013,n1170,kl,q236_1),
       H236_013(h236_013,n1170,kl,q237_1),
       H237_013(h237_013,n1170,kl,q238_1),
       H238_013(h238_013,n1170,kl,q239_1),
       H239_013(h239_013,n1170,kl,q240_1),
       H240_013(h240_013,n1170,kl,q241_1),
       H241_013(h241_013,n1170,kl,q242_1),
       H242_013(h242_013,n1170,kl,q243_1),
       H243_013(h243_013,n1170,kl,q244_1),
       H244_013(h244_013,n1170,kl,q245_1),
       H245_013(h245_013,n1170,kl,q246_1),
       H246_013(h246_013,n1170,kl,q247_1),
       H247_013(h247_013,n1170,kl,q248_1),
       H248_013(h248_013,n1170,kl,q249_1),
       H249_013(h249_013,n1170,kl,q250_1),
       H250_013(h250_013,n1170,kl,q251_1),
       H251_013(h251_013,n1170,kl,q252_1),
       H252_013(h252_013,n1170,kl,q253_1),
       H253_013(h253_013,n1170,kl,q254_1),
       H254_013(h254_013,n1170,kl,q255_1),
       H255_013(h255_013,n1170,kl,q256_1),
       H256_013(h256_013,n1170,kl,q257_1),
       H257_013(h257_013,n1170,kl,q258_1),
       H258_013(h258_013,n1170,kl,q259_1),
       H259_013(h259_013,n1170,kl,q260_1),
       H260_013(h260_013,n1170,kl,q261_1),
       H261_013(h261_013,n1170,kl,q202_1),
       H202_111(h202_111,o1170,q202_0),
       H203_111(h203_111,o1170,q203_0),
       H204_111(h204_111,o1170,q204_0),
       H205_111(h205_111,o1170,q205_0),
       H206_111(h206_111,o1170,q206_0),
       H207_111(h207_111,o1170,q207_0),
       H208_111(h208_111,o1170,q208_0),
       H209_111(h209_111,o1170,q209_0),
       H210_111(h210_111,o1170,q210_0),
       H211_111(h211_111,o1170,q211_0),
       H212_111(h212_111,o1170,q212_0),
       H213_111(h213_111,o1170,q213_0),
       H214_111(h214_111,o1170,q214_0),
       H215_111(h215_111,o1170,q215_0),
       H216_111(h216_111,o1170,q216_0),
       H217_111(h217_111,o1170,q217_0),
       H218_111(h218_111,o1170,q218_0),
       H219_111(h219_111,o1170,q219_0),
       H220_111(h220_111,o1170,q220_0),
       H221_111(h221_111,o1170,q221_0),
       H222_111(h222_111,o1170,q222_0),
       H223_111(h223_111,o1170,q223_0),
       H224_111(h224_111,o1170,q224_0),
       H225_111(h225_111,o1170,q225_0),
       H226_111(h226_111,o1170,q226_0),
       H227_111(h227_111,o1170,q227_0),
       H228_111(h228_111,o1170,q228_0),
       H229_111(h229_111,o1170,q229_0),
       H230_111(h230_111,o1170,q230_0),
       H231_111(h231_111,o1170,q231_0),
       H232_111(h232_111,o1170,q232_0),
       H233_111(h233_111,o1170,q233_0),
       H234_111(h234_111,o1170,q234_0),
       H235_111(h235_111,o1170,q235_0),
       H236_111(h236_111,o1170,q236_0),
       H237_111(h237_111,o1170,q237_0),
       H238_111(h238_111,o1170,q238_0),
       H239_111(h239_111,o1170,q239_0),
       H240_111(h240_111,o1170,q240_0),
       H241_111(h241_111,o1170,q241_0),
       H242_111(h242_111,o1170,q242_0),
       H243_111(h243_111,o1170,q243_0),
       H244_111(h244_111,o1170,q244_0),
       H245_111(h245_111,o1170,q245_0),
       H246_111(h246_111,o1170,q246_0),
       H247_111(h247_111,o1170,q247_0),
       H248_111(h248_111,o1170,q248_0),
       H249_111(h249_111,o1170,q249_0),
       H250_111(h250_111,o1170,q250_0),
       H251_111(h251_111,o1170,q251_0),
       H252_111(h252_111,o1170,q252_0),
       H253_111(h253_111,o1170,q253_0),
       H254_111(h254_111,o1170,q254_0),
       H255_111(h255_111,o1170,q255_0),
       H256_111(h256_111,o1170,q256_0),
       H257_111(h257_111,o1170,q257_0),
       H258_111(h258_111,o1170,q258_0),
       H259_111(h259_111,o1170,q259_0),
       H260_111(h260_111,o1170,q260_0),
       H261_111(h261_111,o1170,q261_0),
       H202_112(h202_112,n1170,q202_1),
       H203_112(h203_112,n1170,q203_1),
       H204_112(h204_112,n1170,q204_1),
       H205_112(h205_112,n1170,q205_1),
       H206_112(h206_112,n1170,q206_1),
       H207_112(h207_112,n1170,q207_1),
       H208_112(h208_112,n1170,q208_1),
       H209_112(h209_112,n1170,q209_1),
       H210_112(h210_112,n1170,q210_1),
       H211_112(h211_112,n1170,q211_1),
       H212_112(h212_112,n1170,q212_1),
       H213_112(h213_112,n1170,q213_1),
       H214_112(h214_112,n1170,q214_1),
       H215_112(h215_112,n1170,q215_1),
       H216_112(h216_112,n1170,q216_1),
       H217_112(h217_112,n1170,q217_1),
       H218_112(h218_112,n1170,q218_1),
       H219_112(h219_112,n1170,q219_1),
       H220_112(h220_112,n1170,q220_1),
       H221_112(h221_112,n1170,q221_1),
       H222_112(h222_112,n1170,q222_1),
       H223_112(h223_112,n1170,q223_1),
       H224_112(h224_112,n1170,q224_1),
       H225_112(h225_112,n1170,q225_1),
       H226_112(h226_112,n1170,q226_1),
       H227_112(h227_112,n1170,q227_1),
       H228_112(h228_112,n1170,q228_1),
       H229_112(h229_112,n1170,q229_1),
       H230_112(h230_112,n1170,q230_1),
       H231_112(h231_112,n1170,q231_1),
       H232_112(h232_112,n1170,q232_1),
       H233_112(h233_112,n1170,q233_1),
       H234_112(h234_112,n1170,q234_1),
       H235_112(h235_112,n1170,q235_1),
       H236_112(h236_112,n1170,q236_1),
       H237_112(h237_112,n1170,q237_1),
       H238_112(h238_112,n1170,q238_1),
       H239_112(h239_112,n1170,q239_1),
       H240_112(h240_112,n1170,q240_1),
       H241_112(h241_112,n1170,q241_1),
       H242_112(h242_112,n1170,q242_1),
       H243_112(h243_112,n1170,q243_1),
       H244_112(h244_112,n1170,q244_1),
       H245_112(h245_112,n1170,q245_1),
       H246_112(h246_112,n1170,q246_1),
       H247_112(h247_112,n1170,q247_1),
       H248_112(h248_112,n1170,q248_1),
       H249_112(h249_112,n1170,q249_1),
       H250_112(h250_112,n1170,q250_1),
       H251_112(h251_112,n1170,q251_1),
       H252_112(h252_112,n1170,q252_1),
       H253_112(h253_112,n1170,q253_1),
       H254_112(h254_112,n1170,q254_1),
       H255_112(h255_112,n1170,q255_1),
       H256_112(h256_112,n1170,q256_1),
       H257_112(h257_112,n1170,q257_1),
       H258_112(h258_112,n1170,q258_1),
       H259_112(h259_112,n1170,q259_1),
       H260_112(h260_112,n1170,q260_1),
       H261_112(h261_112,n1170,q261_1);

or     H00_0(h00_0,h00_011,h00_012),
       H01_0(h01_0,h01_011,h01_012),
       H10_0(h10_0,h10_011,h10_012),
       H11_0(h11_0,h11_011,h11_012),
       H00_1(h00_1,h00_111,h00_112),
       H01_1(h01_1,h01_111,h01_112),
       H10_1(h10_1,h10_111,h10_112),
       H11_1(h11_1,h11_111,h11_112);

and    H00_011(h00_011,o7130,q00_0),
       H01_011(h01_011,o7130,q01_0),
       H10_011(h10_011,o7130,q10_0),
       H11_011(h11_011,o7130,q11_0),
       H00_012(h00_012,n7130,n00_1),
       H01_012(h01_012,n7130,x01_1),
       H10_012(h10_012,n7130,x10_1),
       H11_012(h11_012,n7130,x11_1),
       H00_111(h00_111,o7130,q00_0),
       H01_111(h01_111,o7130,q01_0),
       H10_111(h10_111,o7130,q10_0),
       H11_111(h11_111,o7130,q11_0),
       H00_112(h00_112,n7130,q00_1),
       H01_112(h01_112,n7130,q01_1),
       H10_112(h10_112,n7130,q10_1),
       H11_112(h11_112,n7130,q11_1);

or     Hs_0(hs_0,hs_011,hs_012,n1),
       Hs_1(hs_1,hs_111,hs_112,n1);

and    Hs_011(hs_011,nos,qs_0,o1258),
       Hs_012(hs_012,os,ns_1,o1258),
       Hs_111(hs_111,nos,qs_0,o1258),
       Hs_112(hs_112,os,qs_1,o1258);

or     Hso_0(hso_0,hso_011,hso_012),
       Hso_1(hso_1,hso_111,hso_112);

and    Hso_011(hso_011,o3130,qso_0),
       Hso_012(hso_012,n3130,nso_1),
       Hso_111(hso_111,o3130,qso_0),
       Hso_112(hso_112,n3130,qso_1);

or     H29_0(h29_0,h29_011,h29_012,h29_013,q11_1),
       H30_0(h30_0,h30_011,h30_012,h30_013,q11_1),
       H31_0(h31_0,h31_011,h31_012,h31_013,q11_1),
       H32_0(h32_0,h32_011,h32_012,h32_013,q11_1),
       H33_0(h33_0,h33_011,h33_012,h33_013,q11_1),
       H34_0(h34_0,h34_011,h34_012,h34_013,q11_1),
       H35_0(h35_0,h35_011,h35_012,h35_013,q11_1),
       H36_0(h36_0,h36_011,h36_012,h36_013,q11_1),
       H37_0(h37_0,h37_011,h37_012,h37_013,q11_1),
       H38_0(h38_0,h38_011,h38_012,h38_013,q11_1),
       H39_0(h39_0,h39_011,h39_012,h39_013,q11_1),
       H40_0(h40_0,h40_011,h40_012,h40_013,q11_1),
       H41_0(h41_0,h41_011,h41_012,h41_013,q11_1),
       H42_0(h42_0,h42_011,h42_012,h42_013,q11_1),
       H43_0(h43_0,h43_011,h43_012,h43_013,q11_1),
       H44_0(h44_0,h44_011,h44_012,h44_013),
       H45_0(h45_0,h45_011,h45_012,h45_013),
       H46_0(h46_0,h46_011,h46_012,h46_013),
       H47_0(h47_0,h47_011,h47_012,h47_013),
       H48_0(h48_0,h48_011,h48_012,h48_013),
       H49_0(h49_0,h49_011,h49_012,h49_013),
       H50_0(h50_0,h50_011,h50_012,h50_013),
       H29_1(h29_1,h29_111,h29_112,q11_1),
       H30_1(h30_1,h30_111,h30_112,q11_1),
       H31_1(h31_1,h31_111,h31_112,q11_1),
       H32_1(h32_1,h32_111,h32_112,q11_1),
       H33_1(h33_1,h33_111,h33_112,q11_1),
       H34_1(h34_1,h34_111,h34_112,q11_1),
       H35_1(h35_1,h35_111,h35_112,q11_1),
       H36_1(h36_1,h36_111,h36_112,q11_1),
       H37_1(h37_1,h37_111,h37_112,q11_1),
       H38_1(h38_1,h38_111,h38_112,q11_1),
       H39_1(h39_1,h39_111,h39_112,q11_1),
       H40_1(h40_1,h40_111,h40_112,q11_1),
       H41_1(h41_1,h41_111,h41_112,q11_1),
       H42_1(h42_1,h42_111,h42_112,q11_1),
       H43_1(h43_1,h43_111,h43_112,q11_1),
       H44_1(h44_1,h44_111,h44_112),
       H45_1(h45_1,h45_111,h45_112),
       H46_1(h46_1,h46_111,h46_112),
       H47_1(h47_1,h47_111,h47_112),
       H48_1(h48_1,h48_111,h48_112),
       H49_1(h49_1,h49_111,h49_112),
       H50_1(h50_1,h50_111,h50_112);

and    H29_011(h29_011,nsv,q29_0),
       H30_011(h30_011,nsv,q30_0),
       H31_011(h31_011,nsv,q31_0),
       H32_011(h32_011,nsv,q32_0),
       H33_011(h33_011,nsv,q33_0),
       H34_011(h34_011,nsv,q34_0),
       H35_011(h35_011,nsv,q35_0),
       H36_011(h36_011,nsv,q36_0),
       H37_011(h37_011,nsv,q37_0),
       H38_011(h38_011,nsv,q38_0),
       H39_011(h39_011,nsv,q39_0),
       H40_011(h40_011,nsv,q40_0),
       H41_011(h41_011,nsv,q41_0),
       H42_011(h42_011,nsv,q42_0),
       H43_011(h43_011,nsv,q43_0),
       H44_011(h44_011,nsv,q44_0),
       H45_011(h45_011,nsv,q45_0),
       H46_011(h46_011,nsv,q46_0),
       H47_011(h47_011,nsv,q47_0),
       H48_011(h48_011,nsv,q48_0),
       H49_011(h49_011,nsv,q49_0),
       H50_011(h50_011,nsv,q50_0),
       H29_012(h29_012,asv,sm,dbv1),
       H30_012(h30_012,asv,sm,q29_1),
       H31_012(h31_012,asv,sm,q30_1),
       H32_012(h32_012,asv,sm,q31_1),
       H33_012(h33_012,asv,sm,q32_1),
       H34_012(h34_012,asv,sm,q33_1),
       H35_012(h35_012,asv,sm,q34_1),
       H36_012(h36_012,asv,sm,q35_1),
       H37_012(h37_012,asv,sm,q36_1),
       H38_012(h38_012,asv,sm,q37_1),
       H39_012(h39_012,asv,sm,q38_1),
       H40_012(h40_012,asv,sm,q39_1),
       H41_012(h41_012,asv,sm,q40_1),
       H42_012(h42_012,asv,sm,q41_1),
       H43_012(h43_012,asv,sm,q42_1),
       H44_012(h44_012,asv,sm,q43_1),
       H45_012(h45_012,asv,sm,q44_1),
       H46_012(h46_012,asv,sm,q45_1),
       H47_012(h47_012,asv,sm,q46_1),
       H48_012(h48_012,asv,sm,q47_1),
       H49_012(h49_012,asv,sm,q48_1),
       H50_012(h50_012,asv,sm,q49_1),
       H29_013(h29_013,asv,sp,q30_1),
       H30_013(h30_013,asv,sp,q31_1),
       H31_013(h31_013,asv,sp,q32_1),
       H32_013(h32_013,asv,sp,q33_1),
       H33_013(h33_013,asv,sp,q34_1),
       H34_013(h34_013,asv,sp,q35_1),
       H35_013(h35_013,asv,sp,q36_1),
       H36_013(h36_013,asv,sp,q37_1),
       H37_013(h37_013,asv,sp,q38_1),
       H38_013(h38_013,asv,sp,q39_1),
       H39_013(h39_013,asv,sp,q40_1),
       H40_013(h40_013,asv,sp,q41_1),
       H41_013(h41_013,asv,sp,q42_1),
       H42_013(h42_013,asv,sp,q43_1),
       H43_013(h43_013,asv,sp,q44_1),
       H44_013(h44_013,asv,sp,q45_1),
       H45_013(h45_013,asv,sp,q46_1),
       H46_013(h46_013,asv,sp,q47_1),
       H47_013(h47_013,asv,sp,q48_1),
       H48_013(h48_013,asv,sp,q49_1),
       H49_013(h49_013,asv,sp,q50_1),
       H50_013(h50_013,asv,sp,dbv0),
       H29_111(h29_111,nsv,q29_0),
       H30_111(h30_111,nsv,q30_0),
       H31_111(h31_111,nsv,q31_0),
       H32_111(h32_111,nsv,q32_0),
       H33_111(h33_111,nsv,q33_0),
       H34_111(h34_111,nsv,q34_0),
       H35_111(h35_111,nsv,q35_0),
       H36_111(h36_111,nsv,q36_0),
       H37_111(h37_111,nsv,q37_0),
       H38_111(h38_111,nsv,q38_0),
       H39_111(h39_111,nsv,q39_0),
       H40_111(h40_111,nsv,q40_0),
       H41_111(h41_111,nsv,q41_0),
       H42_111(h42_111,nsv,q42_0),
       H43_111(h43_111,nsv,q43_0),
       H44_111(h44_111,nsv,q44_0),
       H45_111(h45_111,nsv,q45_0),
       H46_111(h46_111,nsv,q46_0),
       H47_111(h47_111,nsv,q47_0),
       H48_111(h48_111,nsv,q48_0),
       H49_111(h49_111,nsv,q49_0),
       H50_111(h50_111,nsv,q50_0),
       H29_112(h29_112,asv,q29_1),
       H30_112(h30_112,asv,q30_1),
       H31_112(h31_112,asv,q31_1),
       H32_112(h32_112,asv,q32_1),
       H33_112(h33_112,asv,q33_1),
       H34_112(h34_112,asv,q34_1),
       H35_112(h35_112,asv,q35_1),
       H36_112(h36_112,asv,q36_1),
       H37_112(h37_112,asv,q37_1),
       H38_112(h38_112,asv,q38_1),
       H39_112(h39_112,asv,q39_1),
       H40_112(h40_112,asv,q40_1),
       H41_112(h41_112,asv,q41_1),
       H42_112(h42_112,asv,q42_1),
       H43_112(h43_112,asv,q43_1),
       H44_112(h44_112,asv,q44_1),
       H45_112(h45_112,asv,q45_1),
       H46_112(h46_112,asv,q46_1),
       H47_112(h47_112,asv,q47_1),
       H48_112(h48_112,asv,q48_1),
       H49_112(h49_112,asv,q49_1),
       H50_112(h50_112,asv,q50_1);

and    Ap102(ap102,q102_1,q000010_1),
       Ap103(ap103,q103_1,q000011_1),
       Ap104(ap104,q104_1,q000100_1),
       Ap105(ap105,q105_1,q000101_1),
       Ap106(ap106,q106_1,q000110_1),
       Ap107(ap107,q107_1,q000111_1),
       Ap108(ap108,q108_1,q001000_1),
       Ap109(ap109,q109_1,q001001_1),
       Ap110(ap110,q110_1,q001010_1),
       Ap111(ap111,q111_1,q001011_1),
       Ap112(ap112,q112_1,q001100_1),
       Ap113(ap113,q113_1,q001101_1),
       Ap114(ap114,q114_1,q001110_1),
       Ap115(ap115,q115_1,q001111_1),
       Ap116(ap116,q116_1,q010000_1),
       Ap117(ap117,q117_1,q010001_1),
       Ap118(ap118,q118_1,q010010_1),
       Ap119(ap119,q119_1,q010011_1),
       Ap120(ap120,q120_1,q010100_1),
       Ap121(ap121,q121_1,q010101_1),
       Ap122(ap122,q122_1,q010110_1),
       Ap123(ap123,q123_1,q010111_1),
       Ap124(ap124,q124_1,q011000_1),
       Ap125(ap125,q125_1,q011001_1),
       Ap126(ap126,q126_1,q011010_1),
       Ap127(ap127,q127_1,q011011_1),
       Ap128(ap128,q128_1,q011100_1),
       Ap129(ap129,q129_1,q011101_1),
       Ap130(ap130,q130_1,q011110_1),
       Ap131(ap131,q131_1,q011111_1),
       Ap132(ap132,q132_1,q100000_1),
       Ap133(ap133,q133_1,q100001_1),
       Ap134(ap134,q134_1,q100010_1),
       Ap135(ap135,q135_1,q100011_1),
       Ap136(ap136,q136_1,q100100_1),
       Ap137(ap137,q137_1,q100101_1),
       Ap138(ap138,q138_1,q100110_1),
       Ap139(ap139,q139_1,q100111_1),
       Ap140(ap140,q140_1,q101000_1),
       Ap141(ap141,q141_1,q101001_1),
       Ap142(ap142,q142_1,q101010_1),
       Ap143(ap143,q143_1,q101011_1),
       Ap144(ap144,q144_1,q101100_1),
       Ap145(ap145,q145_1,q101101_1),
       Ap146(ap146,q146_1,q101110_1),
       Ap147(ap147,q147_1,q101111_1),
       Ap148(ap148,q148_1,q110000_1),
       Ap149(ap149,q149_1,q110001_1),
       Ap150(ap150,q150_1,q110010_1),
       Ap151(ap151,q151_1,q110011_1),
       Ap152(ap152,q152_1,q110100_1),
       Ap153(ap153,q153_1,q110101_1),
       Ap154(ap154,q154_1,q110110_1),
       Ap155(ap155,q155_1,q110111_1),
       Ap156(ap156,q156_1,q111000_1),
       Ap157(ap157,q157_1,q111001_1),
       Ap158(ap158,q158_1,q111010_1),
       Ap159(ap159,q159_1,q111011_1),
       Ap160(ap160,q160_1,q111100_1),
       Ap161(ap161,q161_1,q111101_1),
       Ap202(ap202,q202_1,q000010_1),
       Ap203(ap203,q203_1,q000011_1),
       Ap204(ap204,q204_1,q000100_1),
       Ap205(ap205,q205_1,q000101_1),
       Ap206(ap206,q206_1,q000110_1),
       Ap207(ap207,q207_1,q000111_1),
       Ap208(ap208,q208_1,q001000_1),
       Ap209(ap209,q209_1,q001001_1),
       Ap210(ap210,q210_1,q001010_1),
       Ap211(ap211,q211_1,q001011_1),
       Ap212(ap212,q212_1,q001100_1),
       Ap213(ap213,q213_1,q001101_1),
       Ap214(ap214,q214_1,q001110_1),
       Ap215(ap215,q215_1,q001111_1),
       Ap216(ap216,q216_1,q010000_1),
       Ap217(ap217,q217_1,q010001_1),
       Ap218(ap218,q218_1,q010010_1),
       Ap219(ap219,q219_1,q010011_1),
       Ap220(ap220,q220_1,q010100_1),
       Ap221(ap221,q221_1,q010101_1),
       Ap222(ap222,q222_1,q010110_1),
       Ap223(ap223,q223_1,q010111_1),
       Ap224(ap224,q224_1,q011000_1),
       Ap225(ap225,q225_1,q011001_1),
       Ap226(ap226,q226_1,q011010_1),
       Ap227(ap227,q227_1,q011011_1),
       Ap228(ap228,q228_1,q011100_1),
       Ap229(ap229,q229_1,q011101_1),
       Ap230(ap230,q230_1,q011110_1),
       Ap231(ap231,q231_1,q011111_1),
       Ap232(ap232,q232_1,q100000_1),
       Ap233(ap233,q233_1,q100001_1),
       Ap234(ap234,q234_1,q100010_1),
       Ap235(ap235,q235_1,q100011_1),
       Ap236(ap236,q236_1,q100100_1),
       Ap237(ap237,q237_1,q100101_1),
       Ap238(ap238,q238_1,q100110_1),
       Ap239(ap239,q239_1,q100111_1),
       Ap240(ap240,q240_1,q101000_1),
       Ap241(ap241,q241_1,q101001_1),
       Ap242(ap242,q242_1,q101010_1),
       Ap243(ap243,q243_1,q101011_1),
       Ap244(ap244,q244_1,q101100_1),
       Ap245(ap245,q245_1,q101101_1),
       Ap246(ap246,q246_1,q101110_1),
       Ap247(ap247,q247_1,q101111_1),
       Ap248(ap248,q248_1,q110000_1),
       Ap249(ap249,q249_1,q110001_1),
       Ap250(ap250,q250_1,q110010_1),
       Ap251(ap251,q251_1,q110011_1),
       Ap252(ap252,q252_1,q110100_1),
       Ap253(ap253,q253_1,q110101_1),
       Ap254(ap254,q254_1,q110110_1),
       Ap255(ap255,q255_1,q110111_1),
       Ap256(ap256,q256_1,q111000_1),
       Ap257(ap257,q257_1,q111001_1),
       Ap258(ap258,q258_1,q111010_1),
       Ap259(ap259,q259_1,q111011_1),
       Ap260(ap260,q260_1,q111100_1),
       Ap261(ap261,q261_1,q111101_1);

and    Ad10000(ad10000,n163_1,n162_1,n101_1,n100_1),
       Ad10001(ad10001,n163_1,n162_1,n101_1,q100_1),
       Ad10010(ad10010,n163_1,n162_1,q101_1,n100_1),
       Ad10011(ad10011,n163_1,n162_1,q101_1,q100_1),
       Ad10100(ad10100,n163_1,q162_1,n101_1,n100_1),
       Ad10101(ad10101,n163_1,q162_1,n101_1,q100_1),
       Ad10110(ad10110,n163_1,q162_1,q101_1,n100_1),
       Ad10111(ad10111,n163_1,q162_1,q101_1,q100_1),
       Ad11000(ad11000,q163_1,n162_1,n101_1,n100_1),
       Ad11001(ad11001,q163_1,n162_1,n101_1,q100_1),
       Ad11010(ad11010,q163_1,n162_1,q101_1,n100_1),
       Ad11011(ad11011,q163_1,n162_1,q101_1,q100_1),
       Ad11100(ad11100,q163_1,q162_1,n101_1,n100_1),
       Ad11101(ad11101,q163_1,q162_1,n101_1,q100_1),
       Ad11110(ad11110,q163_1,q162_1,q101_1,n100_1),
       Ad11111(ad11111,q163_1,q162_1,q101_1,q100_1),
       Ad20000(ad20000,n263_1,n262_1,n201_1,n200_1),
       Ad20001(ad20001,n263_1,n262_1,n201_1,q200_1),
       Ad20010(ad20010,n263_1,n262_1,q201_1,n200_1),
       Ad20011(ad20011,n263_1,n262_1,q201_1,q200_1),
       Ad20100(ad20100,n263_1,q262_1,n201_1,n200_1),
       Ad20101(ad20101,n263_1,q262_1,n201_1,q200_1),
       Ad20110(ad20110,n263_1,q262_1,q201_1,n200_1),
       Ad20111(ad20111,n263_1,q262_1,q201_1,q200_1),
       Ad21000(ad21000,q263_1,n262_1,n201_1,n200_1),
       Ad21001(ad21001,q263_1,n262_1,n201_1,q200_1),
       Ad21010(ad21010,q263_1,n262_1,q201_1,n200_1),
       Ad21011(ad21011,q263_1,n262_1,q201_1,q200_1),
       Ad21100(ad21100,q263_1,q262_1,n201_1,n200_1),
       Ad21101(ad21101,q263_1,q262_1,n201_1,q200_1),
       Ad21110(ad21110,q263_1,q262_1,q201_1,n200_1),
       Ad21111(ad21111,q263_1,q262_1,q201_1,q200_1);

and    Ams0000(ams0000,n11_1,n10_1,n01_1,n00_1),
       Ams0001(ams0001,n11_1,n10_1,n01_1,q00_1),
       Ams0010(ams0010,n11_1,n10_1,q01_1,n00_1),
       Ams0011(ams0011,n11_1,n10_1,q01_1,q00_1),
       Ams0100(ams0100,n11_1,q10_1,n01_1,n00_1),
       Ams0101(ams0101,n11_1,q10_1,n01_1,q00_1),
       Ams0110(ams0110,n11_1,q10_1,q01_1,n00_1),
       Ams0111(ams0111,n11_1,q10_1,q01_1,q00_1),
       Ams1000(ams1000,q11_1,n10_1,n01_1,n00_1),
       Ams1001(ams1001,q11_1,n10_1,n01_1,q00_1),
       Ams1010(ams1010,q11_1,n10_1,q01_1,n00_1),
       Ams1011(ams1011,q11_1,n10_1,q01_1,q00_1),
       Ams1100(ams1100,q11_1,q10_1,n01_1,n00_1),
       Ams1101(ams1101,q11_1,q10_1,n01_1,q00_1),
       Ams1110(ams1110,q11_1,q10_1,q01_1,n00_1),
       Ams1111(ams1111,q11_1,q10_1,q01_1,q00_1);

not    N100_1(n100_1,q100_1),
       N101_1(n101_1,q101_1),
       N162_1(n162_1,q162_1),
       N163_1(n163_1,q163_1);
xor    X101_1(x101_1,q101_1,q100_1),
       X162_1(x162_1,q162_1,a162_1),
       X163_1(x163_1,q163_1,a163_1);

and    A162_1(a162_1,q101_1,q100_1),
       A163_1(a163_1,a162_1,q162_1);

not    N200_1(n200_1,q200_1),
       N201_1(n201_1,q201_1),
       N262_1(n262_1,q262_1),
       N263_1(n263_1,q263_1);
xor    X201_1(x201_1,q201_1,q200_1),
       X262_1(x262_1,q262_1,a262_1),
       X263_1(x263_1,q263_1,a263_1);

and    A262_1(a262_1,q201_1,q200_1),
       A263_1(a263_1,a262_1,q262_1);

not    N00_1(n00_1,q00_1),
       N01_1(n01_1,q01_1),
       N10_1(n10_1,q10_1),
       N11_1(n11_1,q11_1);
xor    X01_1(x01_1,q01_1,q00_1),
       X10_1(x10_1,q10_1,a10_1),
       X11_1(x11_1,q11_1,a11_1);

and    A10_1(a10_1,q01_1,q00_1),
       A11_1(a11_1,a10_1,q10_1);

or     Od1(od1,ad11010,ad11011,ad11100,ad11101,ad11110,ad11111),
       Od2a(od2a,ad10001,ad10100,ad11011,ad11110),
       Od2b(od2b,ad10101,ad10110,ad11111),
       Od2c(od2c,ad10010,ad11100),
       Od2d(od2d,ad10001,ad10100,ad10111,ad11011,ad11110),
       Od2e(od2e,ad10001,ad10011,ad10100,ad10101,ad10111,ad11001,ad11011,ad11101,ad11110,ad11111),
       Od2f(od2f,ad10001,ad10010,ad10011,ad10111,ad11011,ad11100,ad11101),
       Od2g(od2g,ad10000,ad10001,ad10111,ad11010,ad11011),
       Od3(od3,ad21010,ad21011,ad21100,ad21101,ad21110,ad21111),
       Od4a(od4a,ad20001,ad20100,ad21011,ad21110),
       Od4b(od4b,ad20101,ad20110,ad21111),
       Od4c(od4c,ad20010,ad21100),
       Od4d(od4d,ad20001,ad20100,ad20111,ad21011,ad21110),
       Od4e(od4e,ad20001,ad20011,ad20100,ad20101,ad20111,ad21001,ad21011,ad21101,ad21110,ad21111),
       Od4f(od4f,ad20001,ad20010,ad20011,ad20111,ad21011,ad21100,ad21101),
       Od4g(od4g,ad20000,ad20001,ad20111,ad21010,ad21011);

or     Oms0(oms0,ams1000,ams1010,ams1100),
       Oms1(oms1,ams1110,ams1111),
       Oms(oms,oms0,oms1);

or     Op1(op1,ap102,ap103,ap104,ap105,ap106,ap107,ap108,ap109,ap110,ap111,ap112,ap113,ap114,ap115,ap116,ap117,ap118,ap119,ap120,ap121,ap122,ap123,ap124,ap125,ap126,ap127,ap128,ap129,ap130,ap131,ap132,ap133,ap134,ap135,ap136,ap137,ap138,ap139,ap140,ap141,ap142,ap143,ap144,ap145,ap146,ap147,ap148,ap149,ap150,ap151,ap152,ap153,ap154,ap155,ap156,ap157,ap158,ap159,ap160,ap161),
       Op2(op2,ap202,ap203,ap204,ap205,ap206,ap207,ap208,ap209,ap210,ap211,ap212,ap213,ap214,ap215,ap216,ap217,ap218,ap219,ap220,ap221,ap222,ap223,ap224,ap225,ap226,ap227,ap228,ap229,ap230,ap231,ap232,ap233,ap234,ap235,ap236,ap237,ap238,ap239,ap240,ap241,ap242,ap243,ap244,ap245,ap246,ap247,ap248,ap249,ap250,ap251,ap252,ap253,ap254,ap255,ap256,ap257,ap258,ap259,ap260,ap261);

and    Ap1(ap1,op1,q0000101_1,q0000110_1,q0000111_1),
       Ap2(ap2,op2,q1111010_1,q1111001_1,q1111000_1);

not    N0_0(n0_0,q0_0),
       N1_0(n1_0,q1_0),
       N0000000_1(n0000000_1,q0000000_1),
       N1111111_1(n1111111_1,q1111111_1);

or     H0_0(h0_0,h0_011,h0_012),
       H1_0(h1_0,h1_011,h1_012),
       H0_002(h0_002,ap1,ap2),
       H1_002(h1_002,q000010_1,q111101_1);

and    H0_011(h0_011,h0_021,q0_0),
       H0_012(h0_012,h0_002,q0000101_1,q0000110_1,q0000111_1),
       H1_011(h1_011,h1_021,q1_0),
       H1_012(h1_012,h1_002,q000010_1);

not    H0_021(h0_021,h0_002),
       H1_021(h1_021,h1_002);

not    N1(n1,s1),
       N4(n4,s4),
       N8(n8,s8),
       P1(p1,r1),
       P3(p3,r3);

xor    Xs(xs,sl,sr),
       Xk(xk,kl,kr);

and    Sl(sl,s4,n8),
       Sr(sr,n4,s8),
       Kr(kr,p1,r3),
       Kl(kl,r1,p3);

or     Osv(osv,sp,sm);

and    Asv(asv,osv,h0_002);

not    Nsv(nsv,asv);

xor    X1005(x1005,d5,q163_1),
       X1006(x1006,d6,q162_1),
       X1007(x1007,d7,q101_1),
       X1008(x1008,d8,q100_1),
       X2005(x2005,d5,q263_1),
       X2006(x2006,d6,q262_1),
       X2007(x2007,d7,q201_1),
       X2008(x2008,d8,q200_1);

and    O1258(o1258,o11258,o21258);
or     O11258(o11258,x1005,x1006,x1007,x1008);
or     O21258(o21258,x2005,x2006,x2007,x2008);

or     Os(os,q0000000_1,q1111111_1,aos);

and    Aos(aos,q00_1,q01_1,q10_1,q11_1);

not    Nso_1(nso_1,qso_1);
not    Ns_1(ns_1,qs_1);
not    Nos(nos,os);

or     Sp(sp,sp10,sp11,sp20,sp21),
       Sm(sm,sm10,sm11,sm20,sm21);

and    Sp10(sp10,sr,n1_0,q0000101_1,q0000110_1,q0000111_1),
       Sp11(sp11,sl,q1_0,q0000101_1,q0000110_1,q0000111_1),
       Sp20(sp20,kl,n1_0,q1111010_1,q1111001_1,q1111000_1),
       Sp21(sp21,kr,q1_0,q1111010_1,q1111001_1,q1111000_1),
       Sm10(sm10,sl,n1_0,q0000101_1,q0000110_1,q0000111_1),
       Sm11(sm11,sr,q1_0,q0000101_1,q0000110_1,q0000111_1),
       Sm20(sm20,kr,n1_0,q1111010_1,q1111001_1,q1111000_1),
       Sm21(sm21,kl,q1_0,q1111010_1,q1111001_1,q1111000_1);

not    N0009(n0009,m0009),
       N0010(n0010,m0010),
       N0011(n0011,m0011),
       N0012(n0012,m0012),
       N0013(n0013,m0013),
       N0014(n0014,m0014),
       N0015(n0015,m0015),
       N0016(n0016,m0016),
       N0017(n0017,m0017),
       N0018(n0018,m0018),
       N0019(n0019,m0019);

or     Ld0000(ld0000,m1111111_0,m1111110_0,m1111101_0,m1111100_0,m1111011_0,m1111010_0,m1111001_0,m1111000_0),
       Ld0001(ld0001,m1110111_0,m1110110_0,m1110101_0,m1110100_0,m1110011_0,m1110010_0,m1110001_0,m1110000_0),
       Ld0010(ld0010,m1101111_0,m1101110_0,m1101101_0,m1101100_0,m1101011_0,m1101010_0,m1101001_0,m1101000_0),
       Ld0011(ld0011,m1100111_0,m1100110_0,m1100101_0,m1100100_0,m1100011_0,m1100010_0,m1100001_0,m1100000_0),
       Ld0100(ld0100,m1011111_0,m1011110_0,m1011101_0,m1011100_0,m1011011_0,m1011010_0,m1011001_0,m1011000_0),
       Ld0101(ld0101,m1010111_0,m1010110_0,m1010101_0,m1010100_0,m1010011_0,m1010010_0,m1010001_0,m1010000_0),
       Ld0110(ld0110,m1001111_0,m1001110_0,m1001101_0,m1001100_0,m1001011_0,m1001010_0,m1001001_0,m1001000_0),
       Ld0111(ld0111,m1000111_0,m1000110_0,m1000101_0,m1000100_0,m1000011_0,m1000010_0,m1000001_0,m1000000_0),
       Ld1000(ld1000,m0111111_0,m0111110_0,m0111101_0,m0111100_0,m0111011_0,m0111010_0,m0111001_0,m0111000_0),
       Ld1001(ld1001,m0110111_0,m0110110_0,m0110101_0,m0110100_0,m0110011_0,m0110010_0,m0110001_0,m0110000_0),
       Ld1010(ld1010,m0101111_0,m0101110_0,m0101101_0,m0101100_0,m0101011_0,m0101010_0,m0101001_0,m0101000_0),
       Ld1011(ld1011,m0100111_0,m0100110_0,m0100101_0,m0100100_0,m0100011_0,m0100010_0,m0100001_0,m0100000_0),
       Ld1100(ld1100,m0011111_0,m0011110_0,m0011101_0,m0011100_0,m0011011_0,m0011010_0,m0011001_0,m0011000_0),
       Ld1101(ld1101,m0010111_0,m0010110_0,m0010101_0,m0010100_0,m0010011_0,m0010010_0,m0010001_0,m0010000_0),
       Ld1110(ld1110,m0001111_0,m0001110_0,m0001101_0,m0001100_0,m0001011_0,m0001010_0,m0001001_0,m0001000_0),
       Ld1111(ld1111,m0000111_0,m0000110_0,m0000101_0,m0000100_0,m0000011_0,m0000010_0,m0000001_0,m0000000_0);
/*
assign ld0000=m29_0;
assign ld0001=m30_0;
assign ld0010=m31_0;
assign ld0011=m32_0;
assign ld0100=m33_0;
assign ld0101=m34_0;
assign ld0110=m35_0;
assign ld0111=m36_0;
assign ld1000=m37_0;
assign ld1001=m38_0;
assign ld1010=m39_0;
assign ld1011=m40_0;
assign ld1100=m41_0;
assign ld1101=m42_0;
assign ld1110=m43_0;
assign ld1111=m44_0;
*/
or     G00(l1,m0016,m0015),
       G01(l2,m0016,n0015),
       G10(l3,n0016,m0015),
       G11(l4,n0016,n0015),
       Gup(up,g21,g36,g51,g66),
       Gru(ru,g22,g37,g52,g67),
       Grd(rd,g23,g38,g53,g68),
       Gdn(dn,g24,g39,g54,g69),
       Gld(ld,g25,g40,g55,g70),
       Glu(lu,g26,g41,g56,g71),
       Gml(ml,g27,g42,g57,g72),
       Gmr(mr,g28,g43,g58,g73),
       Gul(ul,g29,g44,g59,g74),
       Gmu(mu,g30,g45,g60,g75),
       Gur(ur,g31,g46,g61,g76),
       Gdl(dl,g32,g47,g62,g77),
       Gmd(md,g33,g48,g63,g78),
       Gdr(dr,g34,g49,g64,g79),
       Gdt(dt,g35,g50,g65,g80);

and    G21(g21,n00,od1),
       G22(g22,n00,dbv0),
       G23(g23,n00,dbv0),
       G24(g24,n00,od1),
       G25(g25,n00,od1),
       G26(g26,n00,od1),
       G27(g27,n00,dbv1),
       G28(g28,n00,dbv1),
       G29(g29,n00,dbv1),
       G30(g30,n00,dbv1),
       G31(g31,n00,dbv1),
       G32(g32,n00,dbv1),
       G33(g33,n00,dbv1),
       G34(g34,n00,dbv1),
       G35(g35,n00,dbv1),
       G36(g36,n01,od2a),
       G37(g37,n01,od2b),
       G38(g38,n01,od2c),
       G39(g39,n01,od2d),
       G40(g40,n01,od2e),
       G41(g41,n01,od2f),
       G42(g42,n01,od2g),
       G43(g43,n01,od2g),
       G44(g44,n01,dbv1),
       G45(g45,n01,dbv1),
       G46(g46,n01,dbv1),
       G47(g47,n01,dbv1),
       G48(g48,n01,dbv1),
       G49(g49,n01,dbv1),
       G50(g50,n01,dbv1),
       G51(g51,n10,od3),
       G52(g52,n10,dbv0),
       G53(g53,n10,dbv0),
       G54(g54,n10,od3),
       G55(g55,n10,od3),
       G56(g56,n10,od3),
       G57(g57,n10,dbv1),
       G58(g58,n10,dbv1),
       G59(g59,n10,dbv1),
       G60(g60,n10,dbv1),
       G61(g61,n10,dbv1),
       G62(g62,n10,dbv1),
       G63(g63,n10,dbv1),
       G64(g64,n10,dbv1),
       G65(g65,n10,dbv1),
       G66(g66,n11,od4a),
       G67(g67,n11,od4b),
       G68(g68,n11,od4c),
       G69(g69,n11,od4d),
       G70(g70,n11,od4e),
       G71(g71,n11,od4f),
       G72(g72,n11,od4g),
       G73(g73,n11,od4g),
       G74(g74,n11,dbv1),
       G75(g75,n11,dbv1),
       G76(g76,n11,dbv1),
       G77(g77,n11,dbv1),
       G78(g78,n11,dbv1),
       G79(g79,n11,dbv1),
       G80(g80,n11,dbv1);

not    N00(n00,l1),
       N01(n01,l2),
       N10(n10,l3),
       N11(n11,l4);

assign c4=0;

assign appsel=1;
assign bck=m0333;
assign data=xdata;
assign sysclk=clk;
assign ws=m0338;

xor    Xdata(xdata,adata,mso_0);
and    Adata(adata,m0336,m0335,m0334);

assign cs1=n0016;
assign cs2=m0016;
assign dbv0=0;
assign dbv1=1;
assign di=m0011;
assign en=m0008;
assign rst=1;
assign rw=0;

or     Db0(db0,adb000,adb001,adb010,adb011,adb00000000000,adb00000000001,adb00000000010,adb00000000011,adb00000000100,adb00000000101,adb00000000110,adb00000000111,adb00000001000,adb00000001001,adb00000001010,adb00000001011,adb00000001100,adb00000001101,adb00000001110,adb00000001111,adb00000010000,adb00000010001,adb00000010010,adb00000010011,adb00000010100,adb00000010101,adb00000010110,adb00000010111,adb00000011000,adb00000011001,adb00000011010,adb00000011011,adb00000011100,adb00000011101,adb00000011110,adb00000011111,adb00000100000,adb00000100001,adb00000100010,adb00000100011,adb00000100100,adb00000100101,adb00000100110,adb00000100111,adb00000101000,adb00000101001,adb00000101010,adb00000101011,adb00000101100,adb00000101101,adb00000101110,adb00000101111,adb00000110000,adb00000110001,adb00000110010,adb00000110011,adb00000110100,adb00000110101,adb00000110110,adb00000110111,adb00000111000,adb00000111001,adb00000111010,adb00000111011,adb00000111100,adb00000111101,adb00000111110,adb00000111111,adb00001000000,adb00001000001,adb00001000010,adb00001000011,adb00001000100,adb00001000101,adb00001000110,adb00001000111,adb00001001000,adb00001001001,adb00001001010,adb00001001011,adb00001001100,adb00001001101,adb00001001110,adb00001001111,adb00001010000,adb00001010001,adb00001010010,adb00001010011,adb00001010100,adb00001010101,adb00001010110,adb00001010111,adb00001011000,adb00001011001,adb00001011010,adb00001011011,adb00001011100,adb00001011101,adb00001011110,adb00001011111,adb00001100000,adb00001100001,adb00001100010,adb00001100011,adb00001100100,adb00001100101,adb00001100110,adb00001100111,adb00001101000,adb00001101001,adb00001101010,adb00001101011,adb00001101100,adb00001101101,adb00001101110,adb00001101111,adb00001110000,adb00001110001,adb00001110010,adb00001110011,adb00001110100,adb00001110101,adb00001110110,adb00001110111,adb00001111000,adb00001111001,adb00001111010,adb00001111011,adb00001111100,adb00001111101,adb00001111110,adb00001111111,adb00010000000,adb00010000001,adb00010000010,adb00010000011,adb00010000100,adb00010000101,adb00010000110,adb00010000111,adb00010001000,adb00010001001,adb00010001010,adb00010001011,adb00010001100,adb00010001101,adb00010001110,adb00010001111,adb00010010000,adb00010010001,adb00010010010,adb00010010011,adb00010010100,adb00010010101,adb00010010110,adb00010010111,adb00010011000,adb00010011001,adb00010011010,adb00010011011,adb00010011100,adb00010011101,adb00010011110,adb00010011111,adb00010100000,adb00010100001,adb00010100010,adb00010100011,adb00010100100,adb00010100101,adb00010100110,adb00010100111,adb00010101000,adb00010101001,adb00010101010,adb00010101011,adb00010101100,adb00010101101,adb00010101110,adb00010101111,adb00010110000,adb00010110001,adb00010110010,adb00010110011,adb00010110100,adb00010110101,adb00010110110,adb00010110111,adb00010111000,adb00010111001,adb00010111010,adb00010111011,adb00010111100,adb00010111101,adb00010111110,adb00010111111,adb00011000000,adb00011000001,adb00011000010,adb00011000011,adb00011000100,adb00011000101,adb00011000110,adb00011000111,adb00011001000,adb00011001001,adb00011001010,adb00011001011,adb00011001100,adb00011001101,adb00011001110,adb00011001111,adb00011010000,adb00011010001,adb00011010010,adb00011010011,adb00011010100,adb00011010101,adb00011010110,adb00011010111,adb00011011000,adb00011011001,adb00011011010,adb00011011011,adb00011011100,adb00011011101,adb00011011110,adb00011011111,adb00011100000,adb00011100001,adb00011100010,adb00011100011,adb00011100100,adb00011100101,adb00011100110,adb00011100111,adb00011101000,adb00011101001,adb00011101010,adb00011101011,adb00011101100,adb00011101101,adb00011101110,adb00011101111,adb00011110000,adb00011110001,adb00011110010,adb00011110011,adb00011110100,adb00011110101,adb00011110110,adb00011110111,adb00011111000,adb00011111001,adb00011111010,adb00011111011,adb00011111100,adb00011111101,adb00011111110,adb00011111111,adb00100000000,adb00100000001,adb00100000010,adb00100000011,adb00100000100,adb00100000101,adb00100000110,adb00100000111,adb00100001000,adb00100001001,adb00100001010,adb00100001011,adb00100001100,adb00100001101,adb00100001110,adb00100001111,adb00100010000,adb00100010001,adb00100010010,adb00100010011,adb00100010100,adb00100010101,adb00100010110,adb00100010111,adb00100011000,adb00100011001,adb00100011010,adb00100011011,adb00100011100,adb00100011101,adb00100011110,adb00100011111,adb00100100000,adb00100100001,adb00100100010,adb00100100011,adb00100100100,adb00100100101,adb00100100110,adb00100100111,adb00100101000,adb00100101001,adb00100101010,adb00100101011,adb00100101100,adb00100101101,adb00100101110,adb00100101111,adb00100110000,adb00100110001,adb00100110010,adb00100110011,adb00100110100,adb00100110101,adb00100110110,adb00100110111,adb00100111000,adb00100111001,adb00100111010,adb00100111011,adb00100111100,adb00100111101,adb00100111110,adb00100111111,adb00101000000,adb00101000001,adb00101000010,adb00101000011,adb00101000100,adb00101000101,adb00101000110,adb00101000111,adb00101001000,adb00101001001,adb00101001010,adb00101001011,adb00101001100,adb00101001101,adb00101001110,adb00101001111,adb00101010000,adb00101010001,adb00101010010,adb00101010011,adb00101010100,adb00101010101,adb00101010110,adb00101010111,adb00101011000,adb00101011001,adb00101011010,adb00101011011,adb00101011100,adb00101011101,adb00101011110,adb00101011111,adb00101100000,adb00101100001,adb00101100010,adb00101100011,adb00101100100,adb00101100101,adb00101100110,adb00101100111,adb00101101000,adb00101101001,adb00101101010,adb00101101011,adb00101101100,adb00101101101,adb00101101110,adb00101101111,adb00101110000,adb00101110001,adb00101110010,adb00101110011,adb00101110100,adb00101110101,adb00101110110,adb00101110111,adb00101111000,adb00101111001,adb00101111010,adb00101111011,adb00101111100,adb00101111101,adb00101111110,adb00101111111,adb00110000000,adb00110000001,adb00110000010,adb00110000011,adb00110000100,adb00110000101,adb00110000110,adb00110000111,adb00110001000,adb00110001001,adb00110001010,adb00110001011,adb00110001100,adb00110001101,adb00110001110,adb00110001111,adb00110010000,adb00110010001,adb00110010010,adb00110010011,adb00110010100,adb00110010101,adb00110010110,adb00110010111,adb00110011000,adb00110011001,adb00110011010,adb00110011011,adb00110011100,adb00110011101,adb00110011110,adb00110011111,adb00110100000,adb00110100001,adb00110100010,adb00110100011,adb00110100100,adb00110100101,adb00110100110,adb00110100111,adb00110101000,adb00110101001,adb00110101010,adb00110101011,adb00110101100,adb00110101101,adb00110101110,adb00110101111,adb00110110000,adb00110110001,adb00110110010,adb00110110011,adb00110110100,adb00110110101,adb00110110110,adb00110110111,adb00110111000,adb00110111001,adb00110111010,adb00110111011,adb00110111100,adb00110111101,adb00110111110,adb00110111111,adb00111000000,adb00111000001,adb00111000010,adb00111000011,adb00111000100,adb00111000101,adb00111000110,adb00111000111,adb00111001000,adb00111001001,adb00111001010,adb00111001011,adb00111001100,adb00111001101,adb00111001110,adb00111001111,adb00111010000,adb00111010001,adb00111010010,adb00111010011,adb00111010100,adb00111010101,adb00111010110,adb00111010111,adb00111011000,adb00111011001,adb00111011010,adb00111011011,adb00111011100,adb00111011101,adb00111011110,adb00111011111,adb00111100000,adb00111100001,adb00111100010,adb00111100011,adb00111100100,adb00111100101,adb00111100110,adb00111100111,adb00111101000,adb00111101001,adb00111101010,adb00111101011,adb00111101100,adb00111101101,adb00111101110,adb00111101111,adb00111110000,adb00111110001,adb00111110010,adb00111110011,adb00111110100,adb00111110101,adb00111110110,adb00111110111,adb00111111000,adb00111111001,adb00111111010,adb00111111011,adb00111111100,adb00111111101,adb00111111110,adb00111111111,adb01000000000,adb01000000001,adb01000000010,adb01000000011,adb01000000100,adb01000000101,adb01000000110,adb01000000111,adb01000001000,adb01000001001,adb01000001010,adb01000001011,adb01000001100,adb01000001101,adb01000001110,adb01000001111,adb01000010000,adb01000010001,adb01000010010,adb01000010011,adb01000010100,adb01000010101,adb01000010110,adb01000010111,adb01000011000,adb01000011001,adb01000011010,adb01000011011,adb01000011100,adb01000011101,adb01000011110,adb01000011111,adb01000100000,adb01000100001,adb01000100010,adb01000100011,adb01000100100,adb01000100101,adb01000100110,adb01000100111,adb01000101000,adb01000101001,adb01000101010,adb01000101011,adb01000101100,adb01000101101,adb01000101110,adb01000101111,adb01000110000,adb01000110001,adb01000110010,adb01000110011,adb01000110100,adb01000110101,adb01000110110,adb01000110111,adb01000111000,adb01000111001,adb01000111010,adb01000111011,adb01000111100,adb01000111101,adb01000111110,adb01000111111,adb01001000000,adb01001000001,adb01001000010,adb01001000011,adb01001000100,adb01001000101,adb01001000110,adb01001000111,adb01001001000,adb01001001001,adb01001001010,adb01001001011,adb01001001100,adb01001001101,adb01001001110,adb01001001111,adb01001010000,adb01001010001,adb01001010010,adb01001010011,adb01001010100,adb01001010101,adb01001010110,adb01001010111,adb01001011000,adb01001011001,adb01001011010,adb01001011011,adb01001011100,adb01001011101,adb01001011110,adb01001011111,adb01001100000,adb01001100001,adb01001100010,adb01001100011,adb01001100100,adb01001100101,adb01001100110,adb01001100111,adb01001101000,adb01001101001,adb01001101010,adb01001101011,adb01001101100,adb01001101101,adb01001101110,adb01001101111,adb01001110000,adb01001110001,adb01001110010,adb01001110011,adb01001110100,adb01001110101,adb01001110110,adb01001110111,adb01001111000,adb01001111001,adb01001111010,adb01001111011,adb01001111100,adb01001111101,adb01001111110,adb01001111111,adb01010000000,adb01010000001,adb01010000010,adb01010000011,adb01010000100,adb01010000101,adb01010000110,adb01010000111,adb01010001000,adb01010001001,adb01010001010,adb01010001011,adb01010001100,adb01010001101,adb01010001110,adb01010001111,adb01010010000,adb01010010001,adb01010010010,adb01010010011,adb01010010100,adb01010010101,adb01010010110,adb01010010111,adb01010011000,adb01010011001,adb01010011010,adb01010011011,adb01010011100,adb01010011101,adb01010011110,adb01010011111,adb01010100000,adb01010100001,adb01010100010,adb01010100011,adb01010100100,adb01010100101,adb01010100110,adb01010100111,adb01010101000,adb01010101001,adb01010101010,adb01010101011,adb01010101100,adb01010101101,adb01010101110,adb01010101111,adb01010110000,adb01010110001,adb01010110010,adb01010110011,adb01010110100,adb01010110101,adb01010110110,adb01010110111,adb01010111000,adb01010111001,adb01010111010,adb01010111011,adb01010111100,adb01010111101,adb01010111110,adb01010111111,adb01011000000,adb01011000001,adb01011000010,adb01011000011,adb01011000100,adb01011000101,adb01011000110,adb01011000111,adb01011001000,adb01011001001,adb01011001010,adb01011001011,adb01011001100,adb01011001101,adb01011001110,adb01011001111,adb01011010000,adb01011010001,adb01011010010,adb01011010011,adb01011010100,adb01011010101,adb01011010110,adb01011010111,adb01011011000,adb01011011001,adb01011011010,adb01011011011,adb01011011100,adb01011011101,adb01011011110,adb01011011111,adb01011100000,adb01011100001,adb01011100010,adb01011100011,adb01011100100,adb01011100101,adb01011100110,adb01011100111,adb01011101000,adb01011101001,adb01011101010,adb01011101011,adb01011101100,adb01011101101,adb01011101110,adb01011101111,adb01011110000,adb01011110001,adb01011110010,adb01011110011,adb01011110100,adb01011110101,adb01011110110,adb01011110111,adb01011111000,adb01011111001,adb01011111010,adb01011111011,adb01011111100,adb01011111101,adb01011111110,adb01011111111,adb01100000000,adb01100000001,adb01100000010,adb01100000011,adb01100000100,adb01100000101,adb01100000110,adb01100000111,adb01100001000,adb01100001001,adb01100001010,adb01100001011,adb01100001100,adb01100001101,adb01100001110,adb01100001111,adb01100010000,adb01100010001,adb01100010010,adb01100010011,adb01100010100,adb01100010101,adb01100010110,adb01100010111,adb01100011000,adb01100011001,adb01100011010,adb01100011011,adb01100011100,adb01100011101,adb01100011110,adb01100011111,adb01100100000,adb01100100001,adb01100100010,adb01100100011,adb01100100100,adb01100100101,adb01100100110,adb01100100111,adb01100101000,adb01100101001,adb01100101010,adb01100101011,adb01100101100,adb01100101101,adb01100101110,adb01100101111,adb01100110000,adb01100110001,adb01100110010,adb01100110011,adb01100110100,adb01100110101,adb01100110110,adb01100110111,adb01100111000,adb01100111001,adb01100111010,adb01100111011,adb01100111100,adb01100111101,adb01100111110,adb01100111111,adb01101000000,adb01101000001,adb01101000010,adb01101000011,adb01101000100,adb01101000101,adb01101000110,adb01101000111,adb01101001000,adb01101001001,adb01101001010,adb01101001011,adb01101001100,adb01101001101,adb01101001110,adb01101001111,adb01101010000,adb01101010001,adb01101010010,adb01101010011,adb01101010100,adb01101010101,adb01101010110,adb01101010111,adb01101011000,adb01101011001,adb01101011010,adb01101011011,adb01101011100,adb01101011101,adb01101011110,adb01101011111,adb01101100000,adb01101100001,adb01101100010,adb01101100011,adb01101100100,adb01101100101,adb01101100110,adb01101100111,adb01101101000,adb01101101001,adb01101101010,adb01101101011,adb01101101100,adb01101101101,adb01101101110,adb01101101111,adb01101110000,adb01101110001,adb01101110010,adb01101110011,adb01101110100,adb01101110101,adb01101110110,adb01101110111,adb01101111000,adb01101111001,adb01101111010,adb01101111011,adb01101111100,adb01101111101,adb01101111110,adb01101111111,adb01110000000,adb01110000001,adb01110000010,adb01110000011,adb01110000100,adb01110000101,adb01110000110,adb01110000111,adb01110001000,adb01110001001,adb01110001010,adb01110001011,adb01110001100,adb01110001101,adb01110001110,adb01110001111,adb01110010000,adb01110010001,adb01110010010,adb01110010011,adb01110010100,adb01110010101,adb01110010110,adb01110010111,adb01110011000,adb01110011001,adb01110011010,adb01110011011,adb01110011100,adb01110011101,adb01110011110,adb01110011111,adb01110100000,adb01110100001,adb01110100010,adb01110100011,adb01110100100,adb01110100101,adb01110100110,adb01110100111,adb01110101000,adb01110101001,adb01110101010,adb01110101011,adb01110101100,adb01110101101,adb01110101110,adb01110101111,adb01110110000,adb01110110001,adb01110110010,adb01110110011,adb01110110100,adb01110110101,adb01110110110,adb01110110111,adb01110111000,adb01110111001,adb01110111010,adb01110111011,adb01110111100,adb01110111101,adb01110111110,adb01110111111,adb01111000000,adb01111000001,adb01111000010,adb01111000011,adb01111000100,adb01111000101,adb01111000110,adb01111000111,adb01111001000,adb01111001001,adb01111001010,adb01111001011,adb01111001100,adb01111001101,adb01111001110,adb01111001111,adb01111010000,adb01111010001,adb01111010010,adb01111010011,adb01111010100,adb01111010101,adb01111010110,adb01111010111,adb01111011000,adb01111011001,adb01111011010,adb01111011011,adb01111011100,adb01111011101,adb01111011110,adb01111011111,adb01111100000,adb01111100001,adb01111100010,adb01111100011,adb01111100100,adb01111100101,adb01111100110,adb01111100111,adb01111101000,adb01111101001,adb01111101010,adb01111101011,adb01111101100,adb01111101101,adb01111101110,adb01111101111,adb01111110000,adb01111110001,adb01111110010,adb01111110011,adb01111110100,adb01111110101,adb01111110110,adb01111110111,adb01111111000,adb01111111001,adb01111111010,adb01111111011,adb01111111100,adb01111111101,adb01111111110,adb01111111111,adbp107,adbp115,adbp123,adbp131,adbp139,adbp147,adbp155,adbp207,adbp215,adbp223,adbp231,adbp239,adbp247,adbp255,adbtopline0),
       Db1(db1,adb100,adb101,adb110,adb111,adb10000000000,adb10000000001,adb10000000010,adb10000000011,adb10000000100,adb10000000101,adb10000000110,adb10000000111,adb10000001000,adb10000001001,adb10000001010,adb10000001011,adb10000001100,adb10000001101,adb10000001110,adb10000001111,adb10000010000,adb10000010001,adb10000010010,adb10000010011,adb10000010100,adb10000010101,adb10000010110,adb10000010111,adb10000011000,adb10000011001,adb10000011010,adb10000011011,adb10000011100,adb10000011101,adb10000011110,adb10000011111,adb10000100000,adb10000100001,adb10000100010,adb10000100011,adb10000100100,adb10000100101,adb10000100110,adb10000100111,adb10000101000,adb10000101001,adb10000101010,adb10000101011,adb10000101100,adb10000101101,adb10000101110,adb10000101111,adb10000110000,adb10000110001,adb10000110010,adb10000110011,adb10000110100,adb10000110101,adb10000110110,adb10000110111,adb10000111000,adb10000111001,adb10000111010,adb10000111011,adb10000111100,adb10000111101,adb10000111110,adb10000111111,adb10001000000,adb10001000001,adb10001000010,adb10001000011,adb10001000100,adb10001000101,adb10001000110,adb10001000111,adb10001001000,adb10001001001,adb10001001010,adb10001001011,adb10001001100,adb10001001101,adb10001001110,adb10001001111,adb10001010000,adb10001010001,adb10001010010,adb10001010011,adb10001010100,adb10001010101,adb10001010110,adb10001010111,adb10001011000,adb10001011001,adb10001011010,adb10001011011,adb10001011100,adb10001011101,adb10001011110,adb10001011111,adb10001100000,adb10001100001,adb10001100010,adb10001100011,adb10001100100,adb10001100101,adb10001100110,adb10001100111,adb10001101000,adb10001101001,adb10001101010,adb10001101011,adb10001101100,adb10001101101,adb10001101110,adb10001101111,adb10001110000,adb10001110001,adb10001110010,adb10001110011,adb10001110100,adb10001110101,adb10001110110,adb10001110111,adb10001111000,adb10001111001,adb10001111010,adb10001111011,adb10001111100,adb10001111101,adb10001111110,adb10001111111,adb10010000000,adb10010000001,adb10010000010,adb10010000011,adb10010000100,adb10010000101,adb10010000110,adb10010000111,adb10010001000,adb10010001001,adb10010001010,adb10010001011,adb10010001100,adb10010001101,adb10010001110,adb10010001111,adb10010010000,adb10010010001,adb10010010010,adb10010010011,adb10010010100,adb10010010101,adb10010010110,adb10010010111,adb10010011000,adb10010011001,adb10010011010,adb10010011011,adb10010011100,adb10010011101,adb10010011110,adb10010011111,adb10010100000,adb10010100001,adb10010100010,adb10010100011,adb10010100100,adb10010100101,adb10010100110,adb10010100111,adb10010101000,adb10010101001,adb10010101010,adb10010101011,adb10010101100,adb10010101101,adb10010101110,adb10010101111,adb10010110000,adb10010110001,adb10010110010,adb10010110011,adb10010110100,adb10010110101,adb10010110110,adb10010110111,adb10010111000,adb10010111001,adb10010111010,adb10010111011,adb10010111100,adb10010111101,adb10010111110,adb10010111111,adb10011000000,adb10011000001,adb10011000010,adb10011000011,adb10011000100,adb10011000101,adb10011000110,adb10011000111,adb10011001000,adb10011001001,adb10011001010,adb10011001011,adb10011001100,adb10011001101,adb10011001110,adb10011001111,adb10011010000,adb10011010001,adb10011010010,adb10011010011,adb10011010100,adb10011010101,adb10011010110,adb10011010111,adb10011011000,adb10011011001,adb10011011010,adb10011011011,adb10011011100,adb10011011101,adb10011011110,adb10011011111,adb10011100000,adb10011100001,adb10011100010,adb10011100011,adb10011100100,adb10011100101,adb10011100110,adb10011100111,adb10011101000,adb10011101001,adb10011101010,adb10011101011,adb10011101100,adb10011101101,adb10011101110,adb10011101111,adb10011110000,adb10011110001,adb10011110010,adb10011110011,adb10011110100,adb10011110101,adb10011110110,adb10011110111,adb10011111000,adb10011111001,adb10011111010,adb10011111011,adb10011111100,adb10011111101,adb10011111110,adb10011111111,adb10100000000,adb10100000001,adb10100000010,adb10100000011,adb10100000100,adb10100000101,adb10100000110,adb10100000111,adb10100001000,adb10100001001,adb10100001010,adb10100001011,adb10100001100,adb10100001101,adb10100001110,adb10100001111,adb10100010000,adb10100010001,adb10100010010,adb10100010011,adb10100010100,adb10100010101,adb10100010110,adb10100010111,adb10100011000,adb10100011001,adb10100011010,adb10100011011,adb10100011100,adb10100011101,adb10100011110,adb10100011111,adb10100100000,adb10100100001,adb10100100010,adb10100100011,adb10100100100,adb10100100101,adb10100100110,adb10100100111,adb10100101000,adb10100101001,adb10100101010,adb10100101011,adb10100101100,adb10100101101,adb10100101110,adb10100101111,adb10100110000,adb10100110001,adb10100110010,adb10100110011,adb10100110100,adb10100110101,adb10100110110,adb10100110111,adb10100111000,adb10100111001,adb10100111010,adb10100111011,adb10100111100,adb10100111101,adb10100111110,adb10100111111,adb10101000000,adb10101000001,adb10101000010,adb10101000011,adb10101000100,adb10101000101,adb10101000110,adb10101000111,adb10101001000,adb10101001001,adb10101001010,adb10101001011,adb10101001100,adb10101001101,adb10101001110,adb10101001111,adb10101010000,adb10101010001,adb10101010010,adb10101010011,adb10101010100,adb10101010101,adb10101010110,adb10101010111,adb10101011000,adb10101011001,adb10101011010,adb10101011011,adb10101011100,adb10101011101,adb10101011110,adb10101011111,adb10101100000,adb10101100001,adb10101100010,adb10101100011,adb10101100100,adb10101100101,adb10101100110,adb10101100111,adb10101101000,adb10101101001,adb10101101010,adb10101101011,adb10101101100,adb10101101101,adb10101101110,adb10101101111,adb10101110000,adb10101110001,adb10101110010,adb10101110011,adb10101110100,adb10101110101,adb10101110110,adb10101110111,adb10101111000,adb10101111001,adb10101111010,adb10101111011,adb10101111100,adb10101111101,adb10101111110,adb10101111111,adb10110000000,adb10110000001,adb10110000010,adb10110000011,adb10110000100,adb10110000101,adb10110000110,adb10110000111,adb10110001000,adb10110001001,adb10110001010,adb10110001011,adb10110001100,adb10110001101,adb10110001110,adb10110001111,adb10110010000,adb10110010001,adb10110010010,adb10110010011,adb10110010100,adb10110010101,adb10110010110,adb10110010111,adb10110011000,adb10110011001,adb10110011010,adb10110011011,adb10110011100,adb10110011101,adb10110011110,adb10110011111,adb10110100000,adb10110100001,adb10110100010,adb10110100011,adb10110100100,adb10110100101,adb10110100110,adb10110100111,adb10110101000,adb10110101001,adb10110101010,adb10110101011,adb10110101100,adb10110101101,adb10110101110,adb10110101111,adb10110110000,adb10110110001,adb10110110010,adb10110110011,adb10110110100,adb10110110101,adb10110110110,adb10110110111,adb10110111000,adb10110111001,adb10110111010,adb10110111011,adb10110111100,adb10110111101,adb10110111110,adb10110111111,adb10111000000,adb10111000001,adb10111000010,adb10111000011,adb10111000100,adb10111000101,adb10111000110,adb10111000111,adb10111001000,adb10111001001,adb10111001010,adb10111001011,adb10111001100,adb10111001101,adb10111001110,adb10111001111,adb10111010000,adb10111010001,adb10111010010,adb10111010011,adb10111010100,adb10111010101,adb10111010110,adb10111010111,adb10111011000,adb10111011001,adb10111011010,adb10111011011,adb10111011100,adb10111011101,adb10111011110,adb10111011111,adb10111100000,adb10111100001,adb10111100010,adb10111100011,adb10111100100,adb10111100101,adb10111100110,adb10111100111,adb10111101000,adb10111101001,adb10111101010,adb10111101011,adb10111101100,adb10111101101,adb10111101110,adb10111101111,adb10111110000,adb10111110001,adb10111110010,adb10111110011,adb10111110100,adb10111110101,adb10111110110,adb10111110111,adb10111111000,adb10111111001,adb10111111010,adb10111111011,adb10111111100,adb10111111101,adb10111111110,adb10111111111,adb11000000000,adb11000000001,adb11000000010,adb11000000011,adb11000000100,adb11000000101,adb11000000110,adb11000000111,adb11000001000,adb11000001001,adb11000001010,adb11000001011,adb11000001100,adb11000001101,adb11000001110,adb11000001111,adb11000010000,adb11000010001,adb11000010010,adb11000010011,adb11000010100,adb11000010101,adb11000010110,adb11000010111,adb11000011000,adb11000011001,adb11000011010,adb11000011011,adb11000011100,adb11000011101,adb11000011110,adb11000011111,adb11000100000,adb11000100001,adb11000100010,adb11000100011,adb11000100100,adb11000100101,adb11000100110,adb11000100111,adb11000101000,adb11000101001,adb11000101010,adb11000101011,adb11000101100,adb11000101101,adb11000101110,adb11000101111,adb11000110000,adb11000110001,adb11000110010,adb11000110011,adb11000110100,adb11000110101,adb11000110110,adb11000110111,adb11000111000,adb11000111001,adb11000111010,adb11000111011,adb11000111100,adb11000111101,adb11000111110,adb11000111111,adb11001000000,adb11001000001,adb11001000010,adb11001000011,adb11001000100,adb11001000101,adb11001000110,adb11001000111,adb11001001000,adb11001001001,adb11001001010,adb11001001011,adb11001001100,adb11001001101,adb11001001110,adb11001001111,adb11001010000,adb11001010001,adb11001010010,adb11001010011,adb11001010100,adb11001010101,adb11001010110,adb11001010111,adb11001011000,adb11001011001,adb11001011010,adb11001011011,adb11001011100,adb11001011101,adb11001011110,adb11001011111,adb11001100000,adb11001100001,adb11001100010,adb11001100011,adb11001100100,adb11001100101,adb11001100110,adb11001100111,adb11001101000,adb11001101001,adb11001101010,adb11001101011,adb11001101100,adb11001101101,adb11001101110,adb11001101111,adb11001110000,adb11001110001,adb11001110010,adb11001110011,adb11001110100,adb11001110101,adb11001110110,adb11001110111,adb11001111000,adb11001111001,adb11001111010,adb11001111011,adb11001111100,adb11001111101,adb11001111110,adb11001111111,adb11010000000,adb11010000001,adb11010000010,adb11010000011,adb11010000100,adb11010000101,adb11010000110,adb11010000111,adb11010001000,adb11010001001,adb11010001010,adb11010001011,adb11010001100,adb11010001101,adb11010001110,adb11010001111,adb11010010000,adb11010010001,adb11010010010,adb11010010011,adb11010010100,adb11010010101,adb11010010110,adb11010010111,adb11010011000,adb11010011001,adb11010011010,adb11010011011,adb11010011100,adb11010011101,adb11010011110,adb11010011111,adb11010100000,adb11010100001,adb11010100010,adb11010100011,adb11010100100,adb11010100101,adb11010100110,adb11010100111,adb11010101000,adb11010101001,adb11010101010,adb11010101011,adb11010101100,adb11010101101,adb11010101110,adb11010101111,adb11010110000,adb11010110001,adb11010110010,adb11010110011,adb11010110100,adb11010110101,adb11010110110,adb11010110111,adb11010111000,adb11010111001,adb11010111010,adb11010111011,adb11010111100,adb11010111101,adb11010111110,adb11010111111,adb11011000000,adb11011000001,adb11011000010,adb11011000011,adb11011000100,adb11011000101,adb11011000110,adb11011000111,adb11011001000,adb11011001001,adb11011001010,adb11011001011,adb11011001100,adb11011001101,adb11011001110,adb11011001111,adb11011010000,adb11011010001,adb11011010010,adb11011010011,adb11011010100,adb11011010101,adb11011010110,adb11011010111,adb11011011000,adb11011011001,adb11011011010,adb11011011011,adb11011011100,adb11011011101,adb11011011110,adb11011011111,adb11011100000,adb11011100001,adb11011100010,adb11011100011,adb11011100100,adb11011100101,adb11011100110,adb11011100111,adb11011101000,adb11011101001,adb11011101010,adb11011101011,adb11011101100,adb11011101101,adb11011101110,adb11011101111,adb11011110000,adb11011110001,adb11011110010,adb11011110011,adb11011110100,adb11011110101,adb11011110110,adb11011110111,adb11011111000,adb11011111001,adb11011111010,adb11011111011,adb11011111100,adb11011111101,adb11011111110,adb11011111111,adb11100000000,adb11100000001,adb11100000010,adb11100000011,adb11100000100,adb11100000101,adb11100000110,adb11100000111,adb11100001000,adb11100001001,adb11100001010,adb11100001011,adb11100001100,adb11100001101,adb11100001110,adb11100001111,adb11100010000,adb11100010001,adb11100010010,adb11100010011,adb11100010100,adb11100010101,adb11100010110,adb11100010111,adb11100011000,adb11100011001,adb11100011010,adb11100011011,adb11100011100,adb11100011101,adb11100011110,adb11100011111,adb11100100000,adb11100100001,adb11100100010,adb11100100011,adb11100100100,adb11100100101,adb11100100110,adb11100100111,adb11100101000,adb11100101001,adb11100101010,adb11100101011,adb11100101100,adb11100101101,adb11100101110,adb11100101111,adb11100110000,adb11100110001,adb11100110010,adb11100110011,adb11100110100,adb11100110101,adb11100110110,adb11100110111,adb11100111000,adb11100111001,adb11100111010,adb11100111011,adb11100111100,adb11100111101,adb11100111110,adb11100111111,adb11101000000,adb11101000001,adb11101000010,adb11101000011,adb11101000100,adb11101000101,adb11101000110,adb11101000111,adb11101001000,adb11101001001,adb11101001010,adb11101001011,adb11101001100,adb11101001101,adb11101001110,adb11101001111,adb11101010000,adb11101010001,adb11101010010,adb11101010011,adb11101010100,adb11101010101,adb11101010110,adb11101010111,adb11101011000,adb11101011001,adb11101011010,adb11101011011,adb11101011100,adb11101011101,adb11101011110,adb11101011111,adb11101100000,adb11101100001,adb11101100010,adb11101100011,adb11101100100,adb11101100101,adb11101100110,adb11101100111,adb11101101000,adb11101101001,adb11101101010,adb11101101011,adb11101101100,adb11101101101,adb11101101110,adb11101101111,adb11101110000,adb11101110001,adb11101110010,adb11101110011,adb11101110100,adb11101110101,adb11101110110,adb11101110111,adb11101111000,adb11101111001,adb11101111010,adb11101111011,adb11101111100,adb11101111101,adb11101111110,adb11101111111,adb11110000000,adb11110000001,adb11110000010,adb11110000011,adb11110000100,adb11110000101,adb11110000110,adb11110000111,adb11110001000,adb11110001001,adb11110001010,adb11110001011,adb11110001100,adb11110001101,adb11110001110,adb11110001111,adb11110010000,adb11110010001,adb11110010010,adb11110010011,adb11110010100,adb11110010101,adb11110010110,adb11110010111,adb11110011000,adb11110011001,adb11110011010,adb11110011011,adb11110011100,adb11110011101,adb11110011110,adb11110011111,adb11110100000,adb11110100001,adb11110100010,adb11110100011,adb11110100100,adb11110100101,adb11110100110,adb11110100111,adb11110101000,adb11110101001,adb11110101010,adb11110101011,adb11110101100,adb11110101101,adb11110101110,adb11110101111,adb11110110000,adb11110110001,adb11110110010,adb11110110011,adb11110110100,adb11110110101,adb11110110110,adb11110110111,adb11110111000,adb11110111001,adb11110111010,adb11110111011,adb11110111100,adb11110111101,adb11110111110,adb11110111111,adb11111000000,adb11111000001,adb11111000010,adb11111000011,adb11111000100,adb11111000101,adb11111000110,adb11111000111,adb11111001000,adb11111001001,adb11111001010,adb11111001011,adb11111001100,adb11111001101,adb11111001110,adb11111001111,adb11111010000,adb11111010001,adb11111010010,adb11111010011,adb11111010100,adb11111010101,adb11111010110,adb11111010111,adb11111011000,adb11111011001,adb11111011010,adb11111011011,adb11111011100,adb11111011101,adb11111011110,adb11111011111,adb11111100000,adb11111100001,adb11111100010,adb11111100011,adb11111100100,adb11111100101,adb11111100110,adb11111100111,adb11111101000,adb11111101001,adb11111101010,adb11111101011,adb11111101100,adb11111101101,adb11111101110,adb11111101111,adb11111110000,adb11111110001,adb11111110010,adb11111110011,adb11111110100,adb11111110101,adb11111110110,adb11111110111,adb11111111000,adb11111111001,adb11111111010,adb11111111011,adb11111111100,adb11111111101,adb11111111110,adb11111111111,adbp106,adbp114,adbp122,adbp130,adbp138,adbp146,adbp154,adbp206,adbp214,adbp222,adbp230,adbp238,adbp246,adbp254,adbtopline0),
       Db2(db2,adb200,adb201,adb210,adb211,adb20000000000,adb20000000001,adb20000000010,adb20000000011,adb20000000100,adb20000000101,adb20000000110,adb20000000111,adb20000001000,adb20000001001,adb20000001010,adb20000001011,adb20000001100,adb20000001101,adb20000001110,adb20000001111,adb20000010000,adb20000010001,adb20000010010,adb20000010011,adb20000010100,adb20000010101,adb20000010110,adb20000010111,adb20000011000,adb20000011001,adb20000011010,adb20000011011,adb20000011100,adb20000011101,adb20000011110,adb20000011111,adb20000100000,adb20000100001,adb20000100010,adb20000100011,adb20000100100,adb20000100101,adb20000100110,adb20000100111,adb20000101000,adb20000101001,adb20000101010,adb20000101011,adb20000101100,adb20000101101,adb20000101110,adb20000101111,adb20000110000,adb20000110001,adb20000110010,adb20000110011,adb20000110100,adb20000110101,adb20000110110,adb20000110111,adb20000111000,adb20000111001,adb20000111010,adb20000111011,adb20000111100,adb20000111101,adb20000111110,adb20000111111,adb20001000000,adb20001000001,adb20001000010,adb20001000011,adb20001000100,adb20001000101,adb20001000110,adb20001000111,adb20001001000,adb20001001001,adb20001001010,adb20001001011,adb20001001100,adb20001001101,adb20001001110,adb20001001111,adb20001010000,adb20001010001,adb20001010010,adb20001010011,adb20001010100,adb20001010101,adb20001010110,adb20001010111,adb20001011000,adb20001011001,adb20001011010,adb20001011011,adb20001011100,adb20001011101,adb20001011110,adb20001011111,adb20001100000,adb20001100001,adb20001100010,adb20001100011,adb20001100100,adb20001100101,adb20001100110,adb20001100111,adb20001101000,adb20001101001,adb20001101010,adb20001101011,adb20001101100,adb20001101101,adb20001101110,adb20001101111,adb20001110000,adb20001110001,adb20001110010,adb20001110011,adb20001110100,adb20001110101,adb20001110110,adb20001110111,adb20001111000,adb20001111001,adb20001111010,adb20001111011,adb20001111100,adb20001111101,adb20001111110,adb20001111111,adb20010000000,adb20010000001,adb20010000010,adb20010000011,adb20010000100,adb20010000101,adb20010000110,adb20010000111,adb20010001000,adb20010001001,adb20010001010,adb20010001011,adb20010001100,adb20010001101,adb20010001110,adb20010001111,adb20010010000,adb20010010001,adb20010010010,adb20010010011,adb20010010100,adb20010010101,adb20010010110,adb20010010111,adb20010011000,adb20010011001,adb20010011010,adb20010011011,adb20010011100,adb20010011101,adb20010011110,adb20010011111,adb20010100000,adb20010100001,adb20010100010,adb20010100011,adb20010100100,adb20010100101,adb20010100110,adb20010100111,adb20010101000,adb20010101001,adb20010101010,adb20010101011,adb20010101100,adb20010101101,adb20010101110,adb20010101111,adb20010110000,adb20010110001,adb20010110010,adb20010110011,adb20010110100,adb20010110101,adb20010110110,adb20010110111,adb20010111000,adb20010111001,adb20010111010,adb20010111011,adb20010111100,adb20010111101,adb20010111110,adb20010111111,adb20011000000,adb20011000001,adb20011000010,adb20011000011,adb20011000100,adb20011000101,adb20011000110,adb20011000111,adb20011001000,adb20011001001,adb20011001010,adb20011001011,adb20011001100,adb20011001101,adb20011001110,adb20011001111,adb20011010000,adb20011010001,adb20011010010,adb20011010011,adb20011010100,adb20011010101,adb20011010110,adb20011010111,adb20011011000,adb20011011001,adb20011011010,adb20011011011,adb20011011100,adb20011011101,adb20011011110,adb20011011111,adb20011100000,adb20011100001,adb20011100010,adb20011100011,adb20011100100,adb20011100101,adb20011100110,adb20011100111,adb20011101000,adb20011101001,adb20011101010,adb20011101011,adb20011101100,adb20011101101,adb20011101110,adb20011101111,adb20011110000,adb20011110001,adb20011110010,adb20011110011,adb20011110100,adb20011110101,adb20011110110,adb20011110111,adb20011111000,adb20011111001,adb20011111010,adb20011111011,adb20011111100,adb20011111101,adb20011111110,adb20011111111,adb20100000000,adb20100000001,adb20100000010,adb20100000011,adb20100000100,adb20100000101,adb20100000110,adb20100000111,adb20100001000,adb20100001001,adb20100001010,adb20100001011,adb20100001100,adb20100001101,adb20100001110,adb20100001111,adb20100010000,adb20100010001,adb20100010010,adb20100010011,adb20100010100,adb20100010101,adb20100010110,adb20100010111,adb20100011000,adb20100011001,adb20100011010,adb20100011011,adb20100011100,adb20100011101,adb20100011110,adb20100011111,adb20100100000,adb20100100001,adb20100100010,adb20100100011,adb20100100100,adb20100100101,adb20100100110,adb20100100111,adb20100101000,adb20100101001,adb20100101010,adb20100101011,adb20100101100,adb20100101101,adb20100101110,adb20100101111,adb20100110000,adb20100110001,adb20100110010,adb20100110011,adb20100110100,adb20100110101,adb20100110110,adb20100110111,adb20100111000,adb20100111001,adb20100111010,adb20100111011,adb20100111100,adb20100111101,adb20100111110,adb20100111111,adb20101000000,adb20101000001,adb20101000010,adb20101000011,adb20101000100,adb20101000101,adb20101000110,adb20101000111,adb20101001000,adb20101001001,adb20101001010,adb20101001011,adb20101001100,adb20101001101,adb20101001110,adb20101001111,adb20101010000,adb20101010001,adb20101010010,adb20101010011,adb20101010100,adb20101010101,adb20101010110,adb20101010111,adb20101011000,adb20101011001,adb20101011010,adb20101011011,adb20101011100,adb20101011101,adb20101011110,adb20101011111,adb20101100000,adb20101100001,adb20101100010,adb20101100011,adb20101100100,adb20101100101,adb20101100110,adb20101100111,adb20101101000,adb20101101001,adb20101101010,adb20101101011,adb20101101100,adb20101101101,adb20101101110,adb20101101111,adb20101110000,adb20101110001,adb20101110010,adb20101110011,adb20101110100,adb20101110101,adb20101110110,adb20101110111,adb20101111000,adb20101111001,adb20101111010,adb20101111011,adb20101111100,adb20101111101,adb20101111110,adb20101111111,adb20110000000,adb20110000001,adb20110000010,adb20110000011,adb20110000100,adb20110000101,adb20110000110,adb20110000111,adb20110001000,adb20110001001,adb20110001010,adb20110001011,adb20110001100,adb20110001101,adb20110001110,adb20110001111,adb20110010000,adb20110010001,adb20110010010,adb20110010011,adb20110010100,adb20110010101,adb20110010110,adb20110010111,adb20110011000,adb20110011001,adb20110011010,adb20110011011,adb20110011100,adb20110011101,adb20110011110,adb20110011111,adb20110100000,adb20110100001,adb20110100010,adb20110100011,adb20110100100,adb20110100101,adb20110100110,adb20110100111,adb20110101000,adb20110101001,adb20110101010,adb20110101011,adb20110101100,adb20110101101,adb20110101110,adb20110101111,adb20110110000,adb20110110001,adb20110110010,adb20110110011,adb20110110100,adb20110110101,adb20110110110,adb20110110111,adb20110111000,adb20110111001,adb20110111010,adb20110111011,adb20110111100,adb20110111101,adb20110111110,adb20110111111,adb20111000000,adb20111000001,adb20111000010,adb20111000011,adb20111000100,adb20111000101,adb20111000110,adb20111000111,adb20111001000,adb20111001001,adb20111001010,adb20111001011,adb20111001100,adb20111001101,adb20111001110,adb20111001111,adb20111010000,adb20111010001,adb20111010010,adb20111010011,adb20111010100,adb20111010101,adb20111010110,adb20111010111,adb20111011000,adb20111011001,adb20111011010,adb20111011011,adb20111011100,adb20111011101,adb20111011110,adb20111011111,adb20111100000,adb20111100001,adb20111100010,adb20111100011,adb20111100100,adb20111100101,adb20111100110,adb20111100111,adb20111101000,adb20111101001,adb20111101010,adb20111101011,adb20111101100,adb20111101101,adb20111101110,adb20111101111,adb20111110000,adb20111110001,adb20111110010,adb20111110011,adb20111110100,adb20111110101,adb20111110110,adb20111110111,adb20111111000,adb20111111001,adb20111111010,adb20111111011,adb20111111100,adb20111111101,adb20111111110,adb20111111111,adb21000000000,adb21000000001,adb21000000010,adb21000000011,adb21000000100,adb21000000101,adb21000000110,adb21000000111,adb21000001000,adb21000001001,adb21000001010,adb21000001011,adb21000001100,adb21000001101,adb21000001110,adb21000001111,adb21000010000,adb21000010001,adb21000010010,adb21000010011,adb21000010100,adb21000010101,adb21000010110,adb21000010111,adb21000011000,adb21000011001,adb21000011010,adb21000011011,adb21000011100,adb21000011101,adb21000011110,adb21000011111,adb21000100000,adb21000100001,adb21000100010,adb21000100011,adb21000100100,adb21000100101,adb21000100110,adb21000100111,adb21000101000,adb21000101001,adb21000101010,adb21000101011,adb21000101100,adb21000101101,adb21000101110,adb21000101111,adb21000110000,adb21000110001,adb21000110010,adb21000110011,adb21000110100,adb21000110101,adb21000110110,adb21000110111,adb21000111000,adb21000111001,adb21000111010,adb21000111011,adb21000111100,adb21000111101,adb21000111110,adb21000111111,adb21001000000,adb21001000001,adb21001000010,adb21001000011,adb21001000100,adb21001000101,adb21001000110,adb21001000111,adb21001001000,adb21001001001,adb21001001010,adb21001001011,adb21001001100,adb21001001101,adb21001001110,adb21001001111,adb21001010000,adb21001010001,adb21001010010,adb21001010011,adb21001010100,adb21001010101,adb21001010110,adb21001010111,adb21001011000,adb21001011001,adb21001011010,adb21001011011,adb21001011100,adb21001011101,adb21001011110,adb21001011111,adb21001100000,adb21001100001,adb21001100010,adb21001100011,adb21001100100,adb21001100101,adb21001100110,adb21001100111,adb21001101000,adb21001101001,adb21001101010,adb21001101011,adb21001101100,adb21001101101,adb21001101110,adb21001101111,adb21001110000,adb21001110001,adb21001110010,adb21001110011,adb21001110100,adb21001110101,adb21001110110,adb21001110111,adb21001111000,adb21001111001,adb21001111010,adb21001111011,adb21001111100,adb21001111101,adb21001111110,adb21001111111,adb21010000000,adb21010000001,adb21010000010,adb21010000011,adb21010000100,adb21010000101,adb21010000110,adb21010000111,adb21010001000,adb21010001001,adb21010001010,adb21010001011,adb21010001100,adb21010001101,adb21010001110,adb21010001111,adb21010010000,adb21010010001,adb21010010010,adb21010010011,adb21010010100,adb21010010101,adb21010010110,adb21010010111,adb21010011000,adb21010011001,adb21010011010,adb21010011011,adb21010011100,adb21010011101,adb21010011110,adb21010011111,adb21010100000,adb21010100001,adb21010100010,adb21010100011,adb21010100100,adb21010100101,adb21010100110,adb21010100111,adb21010101000,adb21010101001,adb21010101010,adb21010101011,adb21010101100,adb21010101101,adb21010101110,adb21010101111,adb21010110000,adb21010110001,adb21010110010,adb21010110011,adb21010110100,adb21010110101,adb21010110110,adb21010110111,adb21010111000,adb21010111001,adb21010111010,adb21010111011,adb21010111100,adb21010111101,adb21010111110,adb21010111111,adb21011000000,adb21011000001,adb21011000010,adb21011000011,adb21011000100,adb21011000101,adb21011000110,adb21011000111,adb21011001000,adb21011001001,adb21011001010,adb21011001011,adb21011001100,adb21011001101,adb21011001110,adb21011001111,adb21011010000,adb21011010001,adb21011010010,adb21011010011,adb21011010100,adb21011010101,adb21011010110,adb21011010111,adb21011011000,adb21011011001,adb21011011010,adb21011011011,adb21011011100,adb21011011101,adb21011011110,adb21011011111,adb21011100000,adb21011100001,adb21011100010,adb21011100011,adb21011100100,adb21011100101,adb21011100110,adb21011100111,adb21011101000,adb21011101001,adb21011101010,adb21011101011,adb21011101100,adb21011101101,adb21011101110,adb21011101111,adb21011110000,adb21011110001,adb21011110010,adb21011110011,adb21011110100,adb21011110101,adb21011110110,adb21011110111,adb21011111000,adb21011111001,adb21011111010,adb21011111011,adb21011111100,adb21011111101,adb21011111110,adb21011111111,adb21100000000,adb21100000001,adb21100000010,adb21100000011,adb21100000100,adb21100000101,adb21100000110,adb21100000111,adb21100001000,adb21100001001,adb21100001010,adb21100001011,adb21100001100,adb21100001101,adb21100001110,adb21100001111,adb21100010000,adb21100010001,adb21100010010,adb21100010011,adb21100010100,adb21100010101,adb21100010110,adb21100010111,adb21100011000,adb21100011001,adb21100011010,adb21100011011,adb21100011100,adb21100011101,adb21100011110,adb21100011111,adb21100100000,adb21100100001,adb21100100010,adb21100100011,adb21100100100,adb21100100101,adb21100100110,adb21100100111,adb21100101000,adb21100101001,adb21100101010,adb21100101011,adb21100101100,adb21100101101,adb21100101110,adb21100101111,adb21100110000,adb21100110001,adb21100110010,adb21100110011,adb21100110100,adb21100110101,adb21100110110,adb21100110111,adb21100111000,adb21100111001,adb21100111010,adb21100111011,adb21100111100,adb21100111101,adb21100111110,adb21100111111,adb21101000000,adb21101000001,adb21101000010,adb21101000011,adb21101000100,adb21101000101,adb21101000110,adb21101000111,adb21101001000,adb21101001001,adb21101001010,adb21101001011,adb21101001100,adb21101001101,adb21101001110,adb21101001111,adb21101010000,adb21101010001,adb21101010010,adb21101010011,adb21101010100,adb21101010101,adb21101010110,adb21101010111,adb21101011000,adb21101011001,adb21101011010,adb21101011011,adb21101011100,adb21101011101,adb21101011110,adb21101011111,adb21101100000,adb21101100001,adb21101100010,adb21101100011,adb21101100100,adb21101100101,adb21101100110,adb21101100111,adb21101101000,adb21101101001,adb21101101010,adb21101101011,adb21101101100,adb21101101101,adb21101101110,adb21101101111,adb21101110000,adb21101110001,adb21101110010,adb21101110011,adb21101110100,adb21101110101,adb21101110110,adb21101110111,adb21101111000,adb21101111001,adb21101111010,adb21101111011,adb21101111100,adb21101111101,adb21101111110,adb21101111111,adb21110000000,adb21110000001,adb21110000010,adb21110000011,adb21110000100,adb21110000101,adb21110000110,adb21110000111,adb21110001000,adb21110001001,adb21110001010,adb21110001011,adb21110001100,adb21110001101,adb21110001110,adb21110001111,adb21110010000,adb21110010001,adb21110010010,adb21110010011,adb21110010100,adb21110010101,adb21110010110,adb21110010111,adb21110011000,adb21110011001,adb21110011010,adb21110011011,adb21110011100,adb21110011101,adb21110011110,adb21110011111,adb21110100000,adb21110100001,adb21110100010,adb21110100011,adb21110100100,adb21110100101,adb21110100110,adb21110100111,adb21110101000,adb21110101001,adb21110101010,adb21110101011,adb21110101100,adb21110101101,adb21110101110,adb21110101111,adb21110110000,adb21110110001,adb21110110010,adb21110110011,adb21110110100,adb21110110101,adb21110110110,adb21110110111,adb21110111000,adb21110111001,adb21110111010,adb21110111011,adb21110111100,adb21110111101,adb21110111110,adb21110111111,adb21111000000,adb21111000001,adb21111000010,adb21111000011,adb21111000100,adb21111000101,adb21111000110,adb21111000111,adb21111001000,adb21111001001,adb21111001010,adb21111001011,adb21111001100,adb21111001101,adb21111001110,adb21111001111,adb21111010000,adb21111010001,adb21111010010,adb21111010011,adb21111010100,adb21111010101,adb21111010110,adb21111010111,adb21111011000,adb21111011001,adb21111011010,adb21111011011,adb21111011100,adb21111011101,adb21111011110,adb21111011111,adb21111100000,adb21111100001,adb21111100010,adb21111100011,adb21111100100,adb21111100101,adb21111100110,adb21111100111,adb21111101000,adb21111101001,adb21111101010,adb21111101011,adb21111101100,adb21111101101,adb21111101110,adb21111101111,adb21111110000,adb21111110001,adb21111110010,adb21111110011,adb21111110100,adb21111110101,adb21111110110,adb21111110111,adb21111111000,adb21111111001,adb21111111010,adb21111111011,adb21111111100,adb21111111101,adb21111111110,adb21111111111,adbp105,adbp113,adbp121,adbp129,adbp137,adbp145,adbp153,adbp161,adbp205,adbp213,adbp221,adbp229,adbp237,adbp245,adbp253,adbp261),
       Db3(db3,adb300,adb301,adb310,adb311,adb30000000000,adb30000000001,adb30000000010,adb30000000011,adb30000000100,adb30000000101,adb30000000110,adb30000000111,adb30000001000,adb30000001001,adb30000001010,adb30000001011,adb30000001100,adb30000001101,adb30000001110,adb30000001111,adb30000010000,adb30000010001,adb30000010010,adb30000010011,adb30000010100,adb30000010101,adb30000010110,adb30000010111,adb30000011000,adb30000011001,adb30000011010,adb30000011011,adb30000011100,adb30000011101,adb30000011110,adb30000011111,adb30000100000,adb30000100001,adb30000100010,adb30000100011,adb30000100100,adb30000100101,adb30000100110,adb30000100111,adb30000101000,adb30000101001,adb30000101010,adb30000101011,adb30000101100,adb30000101101,adb30000101110,adb30000101111,adb30000110000,adb30000110001,adb30000110010,adb30000110011,adb30000110100,adb30000110101,adb30000110110,adb30000110111,adb30000111000,adb30000111001,adb30000111010,adb30000111011,adb30000111100,adb30000111101,adb30000111110,adb30000111111,adb30001000000,adb30001000001,adb30001000010,adb30001000011,adb30001000100,adb30001000101,adb30001000110,adb30001000111,adb30001001000,adb30001001001,adb30001001010,adb30001001011,adb30001001100,adb30001001101,adb30001001110,adb30001001111,adb30001010000,adb30001010001,adb30001010010,adb30001010011,adb30001010100,adb30001010101,adb30001010110,adb30001010111,adb30001011000,adb30001011001,adb30001011010,adb30001011011,adb30001011100,adb30001011101,adb30001011110,adb30001011111,adb30001100000,adb30001100001,adb30001100010,adb30001100011,adb30001100100,adb30001100101,adb30001100110,adb30001100111,adb30001101000,adb30001101001,adb30001101010,adb30001101011,adb30001101100,adb30001101101,adb30001101110,adb30001101111,adb30001110000,adb30001110001,adb30001110010,adb30001110011,adb30001110100,adb30001110101,adb30001110110,adb30001110111,adb30001111000,adb30001111001,adb30001111010,adb30001111011,adb30001111100,adb30001111101,adb30001111110,adb30001111111,adb30010000000,adb30010000001,adb30010000010,adb30010000011,adb30010000100,adb30010000101,adb30010000110,adb30010000111,adb30010001000,adb30010001001,adb30010001010,adb30010001011,adb30010001100,adb30010001101,adb30010001110,adb30010001111,adb30010010000,adb30010010001,adb30010010010,adb30010010011,adb30010010100,adb30010010101,adb30010010110,adb30010010111,adb30010011000,adb30010011001,adb30010011010,adb30010011011,adb30010011100,adb30010011101,adb30010011110,adb30010011111,adb30010100000,adb30010100001,adb30010100010,adb30010100011,adb30010100100,adb30010100101,adb30010100110,adb30010100111,adb30010101000,adb30010101001,adb30010101010,adb30010101011,adb30010101100,adb30010101101,adb30010101110,adb30010101111,adb30010110000,adb30010110001,adb30010110010,adb30010110011,adb30010110100,adb30010110101,adb30010110110,adb30010110111,adb30010111000,adb30010111001,adb30010111010,adb30010111011,adb30010111100,adb30010111101,adb30010111110,adb30010111111,adb30011000000,adb30011000001,adb30011000010,adb30011000011,adb30011000100,adb30011000101,adb30011000110,adb30011000111,adb30011001000,adb30011001001,adb30011001010,adb30011001011,adb30011001100,adb30011001101,adb30011001110,adb30011001111,adb30011010000,adb30011010001,adb30011010010,adb30011010011,adb30011010100,adb30011010101,adb30011010110,adb30011010111,adb30011011000,adb30011011001,adb30011011010,adb30011011011,adb30011011100,adb30011011101,adb30011011110,adb30011011111,adb30011100000,adb30011100001,adb30011100010,adb30011100011,adb30011100100,adb30011100101,adb30011100110,adb30011100111,adb30011101000,adb30011101001,adb30011101010,adb30011101011,adb30011101100,adb30011101101,adb30011101110,adb30011101111,adb30011110000,adb30011110001,adb30011110010,adb30011110011,adb30011110100,adb30011110101,adb30011110110,adb30011110111,adb30011111000,adb30011111001,adb30011111010,adb30011111011,adb30011111100,adb30011111101,adb30011111110,adb30011111111,adb30100000000,adb30100000001,adb30100000010,adb30100000011,adb30100000100,adb30100000101,adb30100000110,adb30100000111,adb30100001000,adb30100001001,adb30100001010,adb30100001011,adb30100001100,adb30100001101,adb30100001110,adb30100001111,adb30100010000,adb30100010001,adb30100010010,adb30100010011,adb30100010100,adb30100010101,adb30100010110,adb30100010111,adb30100011000,adb30100011001,adb30100011010,adb30100011011,adb30100011100,adb30100011101,adb30100011110,adb30100011111,adb30100100000,adb30100100001,adb30100100010,adb30100100011,adb30100100100,adb30100100101,adb30100100110,adb30100100111,adb30100101000,adb30100101001,adb30100101010,adb30100101011,adb30100101100,adb30100101101,adb30100101110,adb30100101111,adb30100110000,adb30100110001,adb30100110010,adb30100110011,adb30100110100,adb30100110101,adb30100110110,adb30100110111,adb30100111000,adb30100111001,adb30100111010,adb30100111011,adb30100111100,adb30100111101,adb30100111110,adb30100111111,adb30101000000,adb30101000001,adb30101000010,adb30101000011,adb30101000100,adb30101000101,adb30101000110,adb30101000111,adb30101001000,adb30101001001,adb30101001010,adb30101001011,adb30101001100,adb30101001101,adb30101001110,adb30101001111,adb30101010000,adb30101010001,adb30101010010,adb30101010011,adb30101010100,adb30101010101,adb30101010110,adb30101010111,adb30101011000,adb30101011001,adb30101011010,adb30101011011,adb30101011100,adb30101011101,adb30101011110,adb30101011111,adb30101100000,adb30101100001,adb30101100010,adb30101100011,adb30101100100,adb30101100101,adb30101100110,adb30101100111,adb30101101000,adb30101101001,adb30101101010,adb30101101011,adb30101101100,adb30101101101,adb30101101110,adb30101101111,adb30101110000,adb30101110001,adb30101110010,adb30101110011,adb30101110100,adb30101110101,adb30101110110,adb30101110111,adb30101111000,adb30101111001,adb30101111010,adb30101111011,adb30101111100,adb30101111101,adb30101111110,adb30101111111,adb30110000000,adb30110000001,adb30110000010,adb30110000011,adb30110000100,adb30110000101,adb30110000110,adb30110000111,adb30110001000,adb30110001001,adb30110001010,adb30110001011,adb30110001100,adb30110001101,adb30110001110,adb30110001111,adb30110010000,adb30110010001,adb30110010010,adb30110010011,adb30110010100,adb30110010101,adb30110010110,adb30110010111,adb30110011000,adb30110011001,adb30110011010,adb30110011011,adb30110011100,adb30110011101,adb30110011110,adb30110011111,adb30110100000,adb30110100001,adb30110100010,adb30110100011,adb30110100100,adb30110100101,adb30110100110,adb30110100111,adb30110101000,adb30110101001,adb30110101010,adb30110101011,adb30110101100,adb30110101101,adb30110101110,adb30110101111,adb30110110000,adb30110110001,adb30110110010,adb30110110011,adb30110110100,adb30110110101,adb30110110110,adb30110110111,adb30110111000,adb30110111001,adb30110111010,adb30110111011,adb30110111100,adb30110111101,adb30110111110,adb30110111111,adb30111000000,adb30111000001,adb30111000010,adb30111000011,adb30111000100,adb30111000101,adb30111000110,adb30111000111,adb30111001000,adb30111001001,adb30111001010,adb30111001011,adb30111001100,adb30111001101,adb30111001110,adb30111001111,adb30111010000,adb30111010001,adb30111010010,adb30111010011,adb30111010100,adb30111010101,adb30111010110,adb30111010111,adb30111011000,adb30111011001,adb30111011010,adb30111011011,adb30111011100,adb30111011101,adb30111011110,adb30111011111,adb30111100000,adb30111100001,adb30111100010,adb30111100011,adb30111100100,adb30111100101,adb30111100110,adb30111100111,adb30111101000,adb30111101001,adb30111101010,adb30111101011,adb30111101100,adb30111101101,adb30111101110,adb30111101111,adb30111110000,adb30111110001,adb30111110010,adb30111110011,adb30111110100,adb30111110101,adb30111110110,adb30111110111,adb30111111000,adb30111111001,adb30111111010,adb30111111011,adb30111111100,adb30111111101,adb30111111110,adb30111111111,adb31000000000,adb31000000001,adb31000000010,adb31000000011,adb31000000100,adb31000000101,adb31000000110,adb31000000111,adb31000001000,adb31000001001,adb31000001010,adb31000001011,adb31000001100,adb31000001101,adb31000001110,adb31000001111,adb31000010000,adb31000010001,adb31000010010,adb31000010011,adb31000010100,adb31000010101,adb31000010110,adb31000010111,adb31000011000,adb31000011001,adb31000011010,adb31000011011,adb31000011100,adb31000011101,adb31000011110,adb31000011111,adb31000100000,adb31000100001,adb31000100010,adb31000100011,adb31000100100,adb31000100101,adb31000100110,adb31000100111,adb31000101000,adb31000101001,adb31000101010,adb31000101011,adb31000101100,adb31000101101,adb31000101110,adb31000101111,adb31000110000,adb31000110001,adb31000110010,adb31000110011,adb31000110100,adb31000110101,adb31000110110,adb31000110111,adb31000111000,adb31000111001,adb31000111010,adb31000111011,adb31000111100,adb31000111101,adb31000111110,adb31000111111,adb31001000000,adb31001000001,adb31001000010,adb31001000011,adb31001000100,adb31001000101,adb31001000110,adb31001000111,adb31001001000,adb31001001001,adb31001001010,adb31001001011,adb31001001100,adb31001001101,adb31001001110,adb31001001111,adb31001010000,adb31001010001,adb31001010010,adb31001010011,adb31001010100,adb31001010101,adb31001010110,adb31001010111,adb31001011000,adb31001011001,adb31001011010,adb31001011011,adb31001011100,adb31001011101,adb31001011110,adb31001011111,adb31001100000,adb31001100001,adb31001100010,adb31001100011,adb31001100100,adb31001100101,adb31001100110,adb31001100111,adb31001101000,adb31001101001,adb31001101010,adb31001101011,adb31001101100,adb31001101101,adb31001101110,adb31001101111,adb31001110000,adb31001110001,adb31001110010,adb31001110011,adb31001110100,adb31001110101,adb31001110110,adb31001110111,adb31001111000,adb31001111001,adb31001111010,adb31001111011,adb31001111100,adb31001111101,adb31001111110,adb31001111111,adb31010000000,adb31010000001,adb31010000010,adb31010000011,adb31010000100,adb31010000101,adb31010000110,adb31010000111,adb31010001000,adb31010001001,adb31010001010,adb31010001011,adb31010001100,adb31010001101,adb31010001110,adb31010001111,adb31010010000,adb31010010001,adb31010010010,adb31010010011,adb31010010100,adb31010010101,adb31010010110,adb31010010111,adb31010011000,adb31010011001,adb31010011010,adb31010011011,adb31010011100,adb31010011101,adb31010011110,adb31010011111,adb31010100000,adb31010100001,adb31010100010,adb31010100011,adb31010100100,adb31010100101,adb31010100110,adb31010100111,adb31010101000,adb31010101001,adb31010101010,adb31010101011,adb31010101100,adb31010101101,adb31010101110,adb31010101111,adb31010110000,adb31010110001,adb31010110010,adb31010110011,adb31010110100,adb31010110101,adb31010110110,adb31010110111,adb31010111000,adb31010111001,adb31010111010,adb31010111011,adb31010111100,adb31010111101,adb31010111110,adb31010111111,adb31011000000,adb31011000001,adb31011000010,adb31011000011,adb31011000100,adb31011000101,adb31011000110,adb31011000111,adb31011001000,adb31011001001,adb31011001010,adb31011001011,adb31011001100,adb31011001101,adb31011001110,adb31011001111,adb31011010000,adb31011010001,adb31011010010,adb31011010011,adb31011010100,adb31011010101,adb31011010110,adb31011010111,adb31011011000,adb31011011001,adb31011011010,adb31011011011,adb31011011100,adb31011011101,adb31011011110,adb31011011111,adb31011100000,adb31011100001,adb31011100010,adb31011100011,adb31011100100,adb31011100101,adb31011100110,adb31011100111,adb31011101000,adb31011101001,adb31011101010,adb31011101011,adb31011101100,adb31011101101,adb31011101110,adb31011101111,adb31011110000,adb31011110001,adb31011110010,adb31011110011,adb31011110100,adb31011110101,adb31011110110,adb31011110111,adb31011111000,adb31011111001,adb31011111010,adb31011111011,adb31011111100,adb31011111101,adb31011111110,adb31011111111,adb31100000000,adb31100000001,adb31100000010,adb31100000011,adb31100000100,adb31100000101,adb31100000110,adb31100000111,adb31100001000,adb31100001001,adb31100001010,adb31100001011,adb31100001100,adb31100001101,adb31100001110,adb31100001111,adb31100010000,adb31100010001,adb31100010010,adb31100010011,adb31100010100,adb31100010101,adb31100010110,adb31100010111,adb31100011000,adb31100011001,adb31100011010,adb31100011011,adb31100011100,adb31100011101,adb31100011110,adb31100011111,adb31100100000,adb31100100001,adb31100100010,adb31100100011,adb31100100100,adb31100100101,adb31100100110,adb31100100111,adb31100101000,adb31100101001,adb31100101010,adb31100101011,adb31100101100,adb31100101101,adb31100101110,adb31100101111,adb31100110000,adb31100110001,adb31100110010,adb31100110011,adb31100110100,adb31100110101,adb31100110110,adb31100110111,adb31100111000,adb31100111001,adb31100111010,adb31100111011,adb31100111100,adb31100111101,adb31100111110,adb31100111111,adb31101000000,adb31101000001,adb31101000010,adb31101000011,adb31101000100,adb31101000101,adb31101000110,adb31101000111,adb31101001000,adb31101001001,adb31101001010,adb31101001011,adb31101001100,adb31101001101,adb31101001110,adb31101001111,adb31101010000,adb31101010001,adb31101010010,adb31101010011,adb31101010100,adb31101010101,adb31101010110,adb31101010111,adb31101011000,adb31101011001,adb31101011010,adb31101011011,adb31101011100,adb31101011101,adb31101011110,adb31101011111,adb31101100000,adb31101100001,adb31101100010,adb31101100011,adb31101100100,adb31101100101,adb31101100110,adb31101100111,adb31101101000,adb31101101001,adb31101101010,adb31101101011,adb31101101100,adb31101101101,adb31101101110,adb31101101111,adb31101110000,adb31101110001,adb31101110010,adb31101110011,adb31101110100,adb31101110101,adb31101110110,adb31101110111,adb31101111000,adb31101111001,adb31101111010,adb31101111011,adb31101111100,adb31101111101,adb31101111110,adb31101111111,adb31110000000,adb31110000001,adb31110000010,adb31110000011,adb31110000100,adb31110000101,adb31110000110,adb31110000111,adb31110001000,adb31110001001,adb31110001010,adb31110001011,adb31110001100,adb31110001101,adb31110001110,adb31110001111,adb31110010000,adb31110010001,adb31110010010,adb31110010011,adb31110010100,adb31110010101,adb31110010110,adb31110010111,adb31110011000,adb31110011001,adb31110011010,adb31110011011,adb31110011100,adb31110011101,adb31110011110,adb31110011111,adb31110100000,adb31110100001,adb31110100010,adb31110100011,adb31110100100,adb31110100101,adb31110100110,adb31110100111,adb31110101000,adb31110101001,adb31110101010,adb31110101011,adb31110101100,adb31110101101,adb31110101110,adb31110101111,adb31110110000,adb31110110001,adb31110110010,adb31110110011,adb31110110100,adb31110110101,adb31110110110,adb31110110111,adb31110111000,adb31110111001,adb31110111010,adb31110111011,adb31110111100,adb31110111101,adb31110111110,adb31110111111,adb31111000000,adb31111000001,adb31111000010,adb31111000011,adb31111000100,adb31111000101,adb31111000110,adb31111000111,adb31111001000,adb31111001001,adb31111001010,adb31111001011,adb31111001100,adb31111001101,adb31111001110,adb31111001111,adb31111010000,adb31111010001,adb31111010010,adb31111010011,adb31111010100,adb31111010101,adb31111010110,adb31111010111,adb31111011000,adb31111011001,adb31111011010,adb31111011011,adb31111011100,adb31111011101,adb31111011110,adb31111011111,adb31111100000,adb31111100001,adb31111100010,adb31111100011,adb31111100100,adb31111100101,adb31111100110,adb31111100111,adb31111101000,adb31111101001,adb31111101010,adb31111101011,adb31111101100,adb31111101101,adb31111101110,adb31111101111,adb31111110000,adb31111110001,adb31111110010,adb31111110011,adb31111110100,adb31111110101,adb31111110110,adb31111110111,adb31111111000,adb31111111001,adb31111111010,adb31111111011,adb31111111100,adb31111111101,adb31111111110,adb31111111111,adbp104,adbp112,adbp120,adbp128,adbp136,adbp144,adbp152,adbp160,adbp204,adbp212,adbp220,adbp228,adbp236,adbp244,adbp252,adbp260),
       Db4(db4,adb400,adb401,adb410,adb411,adb40000000000,adb40000000001,adb40000000010,adb40000000011,adb40000000100,adb40000000101,adb40000000110,adb40000000111,adb40000001000,adb40000001001,adb40000001010,adb40000001011,adb40000001100,adb40000001101,adb40000001110,adb40000001111,adb40000010000,adb40000010001,adb40000010010,adb40000010011,adb40000010100,adb40000010101,adb40000010110,adb40000010111,adb40000011000,adb40000011001,adb40000011010,adb40000011011,adb40000011100,adb40000011101,adb40000011110,adb40000011111,adb40000100000,adb40000100001,adb40000100010,adb40000100011,adb40000100100,adb40000100101,adb40000100110,adb40000100111,adb40000101000,adb40000101001,adb40000101010,adb40000101011,adb40000101100,adb40000101101,adb40000101110,adb40000101111,adb40000110000,adb40000110001,adb40000110010,adb40000110011,adb40000110100,adb40000110101,adb40000110110,adb40000110111,adb40000111000,adb40000111001,adb40000111010,adb40000111011,adb40000111100,adb40000111101,adb40000111110,adb40000111111,adb40001000000,adb40001000001,adb40001000010,adb40001000011,adb40001000100,adb40001000101,adb40001000110,adb40001000111,adb40001001000,adb40001001001,adb40001001010,adb40001001011,adb40001001100,adb40001001101,adb40001001110,adb40001001111,adb40001010000,adb40001010001,adb40001010010,adb40001010011,adb40001010100,adb40001010101,adb40001010110,adb40001010111,adb40001011000,adb40001011001,adb40001011010,adb40001011011,adb40001011100,adb40001011101,adb40001011110,adb40001011111,adb40001100000,adb40001100001,adb40001100010,adb40001100011,adb40001100100,adb40001100101,adb40001100110,adb40001100111,adb40001101000,adb40001101001,adb40001101010,adb40001101011,adb40001101100,adb40001101101,adb40001101110,adb40001101111,adb40001110000,adb40001110001,adb40001110010,adb40001110011,adb40001110100,adb40001110101,adb40001110110,adb40001110111,adb40001111000,adb40001111001,adb40001111010,adb40001111011,adb40001111100,adb40001111101,adb40001111110,adb40001111111,adb40010000000,adb40010000001,adb40010000010,adb40010000011,adb40010000100,adb40010000101,adb40010000110,adb40010000111,adb40010001000,adb40010001001,adb40010001010,adb40010001011,adb40010001100,adb40010001101,adb40010001110,adb40010001111,adb40010010000,adb40010010001,adb40010010010,adb40010010011,adb40010010100,adb40010010101,adb40010010110,adb40010010111,adb40010011000,adb40010011001,adb40010011010,adb40010011011,adb40010011100,adb40010011101,adb40010011110,adb40010011111,adb40010100000,adb40010100001,adb40010100010,adb40010100011,adb40010100100,adb40010100101,adb40010100110,adb40010100111,adb40010101000,adb40010101001,adb40010101010,adb40010101011,adb40010101100,adb40010101101,adb40010101110,adb40010101111,adb40010110000,adb40010110001,adb40010110010,adb40010110011,adb40010110100,adb40010110101,adb40010110110,adb40010110111,adb40010111000,adb40010111001,adb40010111010,adb40010111011,adb40010111100,adb40010111101,adb40010111110,adb40010111111,adb40011000000,adb40011000001,adb40011000010,adb40011000011,adb40011000100,adb40011000101,adb40011000110,adb40011000111,adb40011001000,adb40011001001,adb40011001010,adb40011001011,adb40011001100,adb40011001101,adb40011001110,adb40011001111,adb40011010000,adb40011010001,adb40011010010,adb40011010011,adb40011010100,adb40011010101,adb40011010110,adb40011010111,adb40011011000,adb40011011001,adb40011011010,adb40011011011,adb40011011100,adb40011011101,adb40011011110,adb40011011111,adb40011100000,adb40011100001,adb40011100010,adb40011100011,adb40011100100,adb40011100101,adb40011100110,adb40011100111,adb40011101000,adb40011101001,adb40011101010,adb40011101011,adb40011101100,adb40011101101,adb40011101110,adb40011101111,adb40011110000,adb40011110001,adb40011110010,adb40011110011,adb40011110100,adb40011110101,adb40011110110,adb40011110111,adb40011111000,adb40011111001,adb40011111010,adb40011111011,adb40011111100,adb40011111101,adb40011111110,adb40011111111,adb40100000000,adb40100000001,adb40100000010,adb40100000011,adb40100000100,adb40100000101,adb40100000110,adb40100000111,adb40100001000,adb40100001001,adb40100001010,adb40100001011,adb40100001100,adb40100001101,adb40100001110,adb40100001111,adb40100010000,adb40100010001,adb40100010010,adb40100010011,adb40100010100,adb40100010101,adb40100010110,adb40100010111,adb40100011000,adb40100011001,adb40100011010,adb40100011011,adb40100011100,adb40100011101,adb40100011110,adb40100011111,adb40100100000,adb40100100001,adb40100100010,adb40100100011,adb40100100100,adb40100100101,adb40100100110,adb40100100111,adb40100101000,adb40100101001,adb40100101010,adb40100101011,adb40100101100,adb40100101101,adb40100101110,adb40100101111,adb40100110000,adb40100110001,adb40100110010,adb40100110011,adb40100110100,adb40100110101,adb40100110110,adb40100110111,adb40100111000,adb40100111001,adb40100111010,adb40100111011,adb40100111100,adb40100111101,adb40100111110,adb40100111111,adb40101000000,adb40101000001,adb40101000010,adb40101000011,adb40101000100,adb40101000101,adb40101000110,adb40101000111,adb40101001000,adb40101001001,adb40101001010,adb40101001011,adb40101001100,adb40101001101,adb40101001110,adb40101001111,adb40101010000,adb40101010001,adb40101010010,adb40101010011,adb40101010100,adb40101010101,adb40101010110,adb40101010111,adb40101011000,adb40101011001,adb40101011010,adb40101011011,adb40101011100,adb40101011101,adb40101011110,adb40101011111,adb40101100000,adb40101100001,adb40101100010,adb40101100011,adb40101100100,adb40101100101,adb40101100110,adb40101100111,adb40101101000,adb40101101001,adb40101101010,adb40101101011,adb40101101100,adb40101101101,adb40101101110,adb40101101111,adb40101110000,adb40101110001,adb40101110010,adb40101110011,adb40101110100,adb40101110101,adb40101110110,adb40101110111,adb40101111000,adb40101111001,adb40101111010,adb40101111011,adb40101111100,adb40101111101,adb40101111110,adb40101111111,adb40110000000,adb40110000001,adb40110000010,adb40110000011,adb40110000100,adb40110000101,adb40110000110,adb40110000111,adb40110001000,adb40110001001,adb40110001010,adb40110001011,adb40110001100,adb40110001101,adb40110001110,adb40110001111,adb40110010000,adb40110010001,adb40110010010,adb40110010011,adb40110010100,adb40110010101,adb40110010110,adb40110010111,adb40110011000,adb40110011001,adb40110011010,adb40110011011,adb40110011100,adb40110011101,adb40110011110,adb40110011111,adb40110100000,adb40110100001,adb40110100010,adb40110100011,adb40110100100,adb40110100101,adb40110100110,adb40110100111,adb40110101000,adb40110101001,adb40110101010,adb40110101011,adb40110101100,adb40110101101,adb40110101110,adb40110101111,adb40110110000,adb40110110001,adb40110110010,adb40110110011,adb40110110100,adb40110110101,adb40110110110,adb40110110111,adb40110111000,adb40110111001,adb40110111010,adb40110111011,adb40110111100,adb40110111101,adb40110111110,adb40110111111,adb40111000000,adb40111000001,adb40111000010,adb40111000011,adb40111000100,adb40111000101,adb40111000110,adb40111000111,adb40111001000,adb40111001001,adb40111001010,adb40111001011,adb40111001100,adb40111001101,adb40111001110,adb40111001111,adb40111010000,adb40111010001,adb40111010010,adb40111010011,adb40111010100,adb40111010101,adb40111010110,adb40111010111,adb40111011000,adb40111011001,adb40111011010,adb40111011011,adb40111011100,adb40111011101,adb40111011110,adb40111011111,adb40111100000,adb40111100001,adb40111100010,adb40111100011,adb40111100100,adb40111100101,adb40111100110,adb40111100111,adb40111101000,adb40111101001,adb40111101010,adb40111101011,adb40111101100,adb40111101101,adb40111101110,adb40111101111,adb40111110000,adb40111110001,adb40111110010,adb40111110011,adb40111110100,adb40111110101,adb40111110110,adb40111110111,adb40111111000,adb40111111001,adb40111111010,adb40111111011,adb40111111100,adb40111111101,adb40111111110,adb40111111111,adb41000000000,adb41000000001,adb41000000010,adb41000000011,adb41000000100,adb41000000101,adb41000000110,adb41000000111,adb41000001000,adb41000001001,adb41000001010,adb41000001011,adb41000001100,adb41000001101,adb41000001110,adb41000001111,adb41000010000,adb41000010001,adb41000010010,adb41000010011,adb41000010100,adb41000010101,adb41000010110,adb41000010111,adb41000011000,adb41000011001,adb41000011010,adb41000011011,adb41000011100,adb41000011101,adb41000011110,adb41000011111,adb41000100000,adb41000100001,adb41000100010,adb41000100011,adb41000100100,adb41000100101,adb41000100110,adb41000100111,adb41000101000,adb41000101001,adb41000101010,adb41000101011,adb41000101100,adb41000101101,adb41000101110,adb41000101111,adb41000110000,adb41000110001,adb41000110010,adb41000110011,adb41000110100,adb41000110101,adb41000110110,adb41000110111,adb41000111000,adb41000111001,adb41000111010,adb41000111011,adb41000111100,adb41000111101,adb41000111110,adb41000111111,adb41001000000,adb41001000001,adb41001000010,adb41001000011,adb41001000100,adb41001000101,adb41001000110,adb41001000111,adb41001001000,adb41001001001,adb41001001010,adb41001001011,adb41001001100,adb41001001101,adb41001001110,adb41001001111,adb41001010000,adb41001010001,adb41001010010,adb41001010011,adb41001010100,adb41001010101,adb41001010110,adb41001010111,adb41001011000,adb41001011001,adb41001011010,adb41001011011,adb41001011100,adb41001011101,adb41001011110,adb41001011111,adb41001100000,adb41001100001,adb41001100010,adb41001100011,adb41001100100,adb41001100101,adb41001100110,adb41001100111,adb41001101000,adb41001101001,adb41001101010,adb41001101011,adb41001101100,adb41001101101,adb41001101110,adb41001101111,adb41001110000,adb41001110001,adb41001110010,adb41001110011,adb41001110100,adb41001110101,adb41001110110,adb41001110111,adb41001111000,adb41001111001,adb41001111010,adb41001111011,adb41001111100,adb41001111101,adb41001111110,adb41001111111,adb41010000000,adb41010000001,adb41010000010,adb41010000011,adb41010000100,adb41010000101,adb41010000110,adb41010000111,adb41010001000,adb41010001001,adb41010001010,adb41010001011,adb41010001100,adb41010001101,adb41010001110,adb41010001111,adb41010010000,adb41010010001,adb41010010010,adb41010010011,adb41010010100,adb41010010101,adb41010010110,adb41010010111,adb41010011000,adb41010011001,adb41010011010,adb41010011011,adb41010011100,adb41010011101,adb41010011110,adb41010011111,adb41010100000,adb41010100001,adb41010100010,adb41010100011,adb41010100100,adb41010100101,adb41010100110,adb41010100111,adb41010101000,adb41010101001,adb41010101010,adb41010101011,adb41010101100,adb41010101101,adb41010101110,adb41010101111,adb41010110000,adb41010110001,adb41010110010,adb41010110011,adb41010110100,adb41010110101,adb41010110110,adb41010110111,adb41010111000,adb41010111001,adb41010111010,adb41010111011,adb41010111100,adb41010111101,adb41010111110,adb41010111111,adb41011000000,adb41011000001,adb41011000010,adb41011000011,adb41011000100,adb41011000101,adb41011000110,adb41011000111,adb41011001000,adb41011001001,adb41011001010,adb41011001011,adb41011001100,adb41011001101,adb41011001110,adb41011001111,adb41011010000,adb41011010001,adb41011010010,adb41011010011,adb41011010100,adb41011010101,adb41011010110,adb41011010111,adb41011011000,adb41011011001,adb41011011010,adb41011011011,adb41011011100,adb41011011101,adb41011011110,adb41011011111,adb41011100000,adb41011100001,adb41011100010,adb41011100011,adb41011100100,adb41011100101,adb41011100110,adb41011100111,adb41011101000,adb41011101001,adb41011101010,adb41011101011,adb41011101100,adb41011101101,adb41011101110,adb41011101111,adb41011110000,adb41011110001,adb41011110010,adb41011110011,adb41011110100,adb41011110101,adb41011110110,adb41011110111,adb41011111000,adb41011111001,adb41011111010,adb41011111011,adb41011111100,adb41011111101,adb41011111110,adb41011111111,adb41100000000,adb41100000001,adb41100000010,adb41100000011,adb41100000100,adb41100000101,adb41100000110,adb41100000111,adb41100001000,adb41100001001,adb41100001010,adb41100001011,adb41100001100,adb41100001101,adb41100001110,adb41100001111,adb41100010000,adb41100010001,adb41100010010,adb41100010011,adb41100010100,adb41100010101,adb41100010110,adb41100010111,adb41100011000,adb41100011001,adb41100011010,adb41100011011,adb41100011100,adb41100011101,adb41100011110,adb41100011111,adb41100100000,adb41100100001,adb41100100010,adb41100100011,adb41100100100,adb41100100101,adb41100100110,adb41100100111,adb41100101000,adb41100101001,adb41100101010,adb41100101011,adb41100101100,adb41100101101,adb41100101110,adb41100101111,adb41100110000,adb41100110001,adb41100110010,adb41100110011,adb41100110100,adb41100110101,adb41100110110,adb41100110111,adb41100111000,adb41100111001,adb41100111010,adb41100111011,adb41100111100,adb41100111101,adb41100111110,adb41100111111,adb41101000000,adb41101000001,adb41101000010,adb41101000011,adb41101000100,adb41101000101,adb41101000110,adb41101000111,adb41101001000,adb41101001001,adb41101001010,adb41101001011,adb41101001100,adb41101001101,adb41101001110,adb41101001111,adb41101010000,adb41101010001,adb41101010010,adb41101010011,adb41101010100,adb41101010101,adb41101010110,adb41101010111,adb41101011000,adb41101011001,adb41101011010,adb41101011011,adb41101011100,adb41101011101,adb41101011110,adb41101011111,adb41101100000,adb41101100001,adb41101100010,adb41101100011,adb41101100100,adb41101100101,adb41101100110,adb41101100111,adb41101101000,adb41101101001,adb41101101010,adb41101101011,adb41101101100,adb41101101101,adb41101101110,adb41101101111,adb41101110000,adb41101110001,adb41101110010,adb41101110011,adb41101110100,adb41101110101,adb41101110110,adb41101110111,adb41101111000,adb41101111001,adb41101111010,adb41101111011,adb41101111100,adb41101111101,adb41101111110,adb41101111111,adb41110000000,adb41110000001,adb41110000010,adb41110000011,adb41110000100,adb41110000101,adb41110000110,adb41110000111,adb41110001000,adb41110001001,adb41110001010,adb41110001011,adb41110001100,adb41110001101,adb41110001110,adb41110001111,adb41110010000,adb41110010001,adb41110010010,adb41110010011,adb41110010100,adb41110010101,adb41110010110,adb41110010111,adb41110011000,adb41110011001,adb41110011010,adb41110011011,adb41110011100,adb41110011101,adb41110011110,adb41110011111,adb41110100000,adb41110100001,adb41110100010,adb41110100011,adb41110100100,adb41110100101,adb41110100110,adb41110100111,adb41110101000,adb41110101001,adb41110101010,adb41110101011,adb41110101100,adb41110101101,adb41110101110,adb41110101111,adb41110110000,adb41110110001,adb41110110010,adb41110110011,adb41110110100,adb41110110101,adb41110110110,adb41110110111,adb41110111000,adb41110111001,adb41110111010,adb41110111011,adb41110111100,adb41110111101,adb41110111110,adb41110111111,adb41111000000,adb41111000001,adb41111000010,adb41111000011,adb41111000100,adb41111000101,adb41111000110,adb41111000111,adb41111001000,adb41111001001,adb41111001010,adb41111001011,adb41111001100,adb41111001101,adb41111001110,adb41111001111,adb41111010000,adb41111010001,adb41111010010,adb41111010011,adb41111010100,adb41111010101,adb41111010110,adb41111010111,adb41111011000,adb41111011001,adb41111011010,adb41111011011,adb41111011100,adb41111011101,adb41111011110,adb41111011111,adb41111100000,adb41111100001,adb41111100010,adb41111100011,adb41111100100,adb41111100101,adb41111100110,adb41111100111,adb41111101000,adb41111101001,adb41111101010,adb41111101011,adb41111101100,adb41111101101,adb41111101110,adb41111101111,adb41111110000,adb41111110001,adb41111110010,adb41111110011,adb41111110100,adb41111110101,adb41111110110,adb41111110111,adb41111111000,adb41111111001,adb41111111010,adb41111111011,adb41111111100,adb41111111101,adb41111111110,adb41111111111,adbp103,adbp111,adbp119,adbp127,adbp135,adbp143,adbp151,adbp159,adbp203,adbp211,adbp219,adbp227,adbp235,adbp243,adbp251,adbp259),
       Db5(db5,adb500,adb501,adb510,adb511,adb50000000000,adb50000000001,adb50000000010,adb50000000011,adb50000000100,adb50000000101,adb50000000110,adb50000000111,adb50000001000,adb50000001001,adb50000001010,adb50000001011,adb50000001100,adb50000001101,adb50000001110,adb50000001111,adb50000010000,adb50000010001,adb50000010010,adb50000010011,adb50000010100,adb50000010101,adb50000010110,adb50000010111,adb50000011000,adb50000011001,adb50000011010,adb50000011011,adb50000011100,adb50000011101,adb50000011110,adb50000011111,adb50000100000,adb50000100001,adb50000100010,adb50000100011,adb50000100100,adb50000100101,adb50000100110,adb50000100111,adb50000101000,adb50000101001,adb50000101010,adb50000101011,adb50000101100,adb50000101101,adb50000101110,adb50000101111,adb50000110000,adb50000110001,adb50000110010,adb50000110011,adb50000110100,adb50000110101,adb50000110110,adb50000110111,adb50000111000,adb50000111001,adb50000111010,adb50000111011,adb50000111100,adb50000111101,adb50000111110,adb50000111111,adb50001000000,adb50001000001,adb50001000010,adb50001000011,adb50001000100,adb50001000101,adb50001000110,adb50001000111,adb50001001000,adb50001001001,adb50001001010,adb50001001011,adb50001001100,adb50001001101,adb50001001110,adb50001001111,adb50001010000,adb50001010001,adb50001010010,adb50001010011,adb50001010100,adb50001010101,adb50001010110,adb50001010111,adb50001011000,adb50001011001,adb50001011010,adb50001011011,adb50001011100,adb50001011101,adb50001011110,adb50001011111,adb50001100000,adb50001100001,adb50001100010,adb50001100011,adb50001100100,adb50001100101,adb50001100110,adb50001100111,adb50001101000,adb50001101001,adb50001101010,adb50001101011,adb50001101100,adb50001101101,adb50001101110,adb50001101111,adb50001110000,adb50001110001,adb50001110010,adb50001110011,adb50001110100,adb50001110101,adb50001110110,adb50001110111,adb50001111000,adb50001111001,adb50001111010,adb50001111011,adb50001111100,adb50001111101,adb50001111110,adb50001111111,adb50010000000,adb50010000001,adb50010000010,adb50010000011,adb50010000100,adb50010000101,adb50010000110,adb50010000111,adb50010001000,adb50010001001,adb50010001010,adb50010001011,adb50010001100,adb50010001101,adb50010001110,adb50010001111,adb50010010000,adb50010010001,adb50010010010,adb50010010011,adb50010010100,adb50010010101,adb50010010110,adb50010010111,adb50010011000,adb50010011001,adb50010011010,adb50010011011,adb50010011100,adb50010011101,adb50010011110,adb50010011111,adb50010100000,adb50010100001,adb50010100010,adb50010100011,adb50010100100,adb50010100101,adb50010100110,adb50010100111,adb50010101000,adb50010101001,adb50010101010,adb50010101011,adb50010101100,adb50010101101,adb50010101110,adb50010101111,adb50010110000,adb50010110001,adb50010110010,adb50010110011,adb50010110100,adb50010110101,adb50010110110,adb50010110111,adb50010111000,adb50010111001,adb50010111010,adb50010111011,adb50010111100,adb50010111101,adb50010111110,adb50010111111,adb50011000000,adb50011000001,adb50011000010,adb50011000011,adb50011000100,adb50011000101,adb50011000110,adb50011000111,adb50011001000,adb50011001001,adb50011001010,adb50011001011,adb50011001100,adb50011001101,adb50011001110,adb50011001111,adb50011010000,adb50011010001,adb50011010010,adb50011010011,adb50011010100,adb50011010101,adb50011010110,adb50011010111,adb50011011000,adb50011011001,adb50011011010,adb50011011011,adb50011011100,adb50011011101,adb50011011110,adb50011011111,adb50011100000,adb50011100001,adb50011100010,adb50011100011,adb50011100100,adb50011100101,adb50011100110,adb50011100111,adb50011101000,adb50011101001,adb50011101010,adb50011101011,adb50011101100,adb50011101101,adb50011101110,adb50011101111,adb50011110000,adb50011110001,adb50011110010,adb50011110011,adb50011110100,adb50011110101,adb50011110110,adb50011110111,adb50011111000,adb50011111001,adb50011111010,adb50011111011,adb50011111100,adb50011111101,adb50011111110,adb50011111111,adb50100000000,adb50100000001,adb50100000010,adb50100000011,adb50100000100,adb50100000101,adb50100000110,adb50100000111,adb50100001000,adb50100001001,adb50100001010,adb50100001011,adb50100001100,adb50100001101,adb50100001110,adb50100001111,adb50100010000,adb50100010001,adb50100010010,adb50100010011,adb50100010100,adb50100010101,adb50100010110,adb50100010111,adb50100011000,adb50100011001,adb50100011010,adb50100011011,adb50100011100,adb50100011101,adb50100011110,adb50100011111,adb50100100000,adb50100100001,adb50100100010,adb50100100011,adb50100100100,adb50100100101,adb50100100110,adb50100100111,adb50100101000,adb50100101001,adb50100101010,adb50100101011,adb50100101100,adb50100101101,adb50100101110,adb50100101111,adb50100110000,adb50100110001,adb50100110010,adb50100110011,adb50100110100,adb50100110101,adb50100110110,adb50100110111,adb50100111000,adb50100111001,adb50100111010,adb50100111011,adb50100111100,adb50100111101,adb50100111110,adb50100111111,adb50101000000,adb50101000001,adb50101000010,adb50101000011,adb50101000100,adb50101000101,adb50101000110,adb50101000111,adb50101001000,adb50101001001,adb50101001010,adb50101001011,adb50101001100,adb50101001101,adb50101001110,adb50101001111,adb50101010000,adb50101010001,adb50101010010,adb50101010011,adb50101010100,adb50101010101,adb50101010110,adb50101010111,adb50101011000,adb50101011001,adb50101011010,adb50101011011,adb50101011100,adb50101011101,adb50101011110,adb50101011111,adb50101100000,adb50101100001,adb50101100010,adb50101100011,adb50101100100,adb50101100101,adb50101100110,adb50101100111,adb50101101000,adb50101101001,adb50101101010,adb50101101011,adb50101101100,adb50101101101,adb50101101110,adb50101101111,adb50101110000,adb50101110001,adb50101110010,adb50101110011,adb50101110100,adb50101110101,adb50101110110,adb50101110111,adb50101111000,adb50101111001,adb50101111010,adb50101111011,adb50101111100,adb50101111101,adb50101111110,adb50101111111,adb50110000000,adb50110000001,adb50110000010,adb50110000011,adb50110000100,adb50110000101,adb50110000110,adb50110000111,adb50110001000,adb50110001001,adb50110001010,adb50110001011,adb50110001100,adb50110001101,adb50110001110,adb50110001111,adb50110010000,adb50110010001,adb50110010010,adb50110010011,adb50110010100,adb50110010101,adb50110010110,adb50110010111,adb50110011000,adb50110011001,adb50110011010,adb50110011011,adb50110011100,adb50110011101,adb50110011110,adb50110011111,adb50110100000,adb50110100001,adb50110100010,adb50110100011,adb50110100100,adb50110100101,adb50110100110,adb50110100111,adb50110101000,adb50110101001,adb50110101010,adb50110101011,adb50110101100,adb50110101101,adb50110101110,adb50110101111,adb50110110000,adb50110110001,adb50110110010,adb50110110011,adb50110110100,adb50110110101,adb50110110110,adb50110110111,adb50110111000,adb50110111001,adb50110111010,adb50110111011,adb50110111100,adb50110111101,adb50110111110,adb50110111111,adb50111000000,adb50111000001,adb50111000010,adb50111000011,adb50111000100,adb50111000101,adb50111000110,adb50111000111,adb50111001000,adb50111001001,adb50111001010,adb50111001011,adb50111001100,adb50111001101,adb50111001110,adb50111001111,adb50111010000,adb50111010001,adb50111010010,adb50111010011,adb50111010100,adb50111010101,adb50111010110,adb50111010111,adb50111011000,adb50111011001,adb50111011010,adb50111011011,adb50111011100,adb50111011101,adb50111011110,adb50111011111,adb50111100000,adb50111100001,adb50111100010,adb50111100011,adb50111100100,adb50111100101,adb50111100110,adb50111100111,adb50111101000,adb50111101001,adb50111101010,adb50111101011,adb50111101100,adb50111101101,adb50111101110,adb50111101111,adb50111110000,adb50111110001,adb50111110010,adb50111110011,adb50111110100,adb50111110101,adb50111110110,adb50111110111,adb50111111000,adb50111111001,adb50111111010,adb50111111011,adb50111111100,adb50111111101,adb50111111110,adb50111111111,adb51000000000,adb51000000001,adb51000000010,adb51000000011,adb51000000100,adb51000000101,adb51000000110,adb51000000111,adb51000001000,adb51000001001,adb51000001010,adb51000001011,adb51000001100,adb51000001101,adb51000001110,adb51000001111,adb51000010000,adb51000010001,adb51000010010,adb51000010011,adb51000010100,adb51000010101,adb51000010110,adb51000010111,adb51000011000,adb51000011001,adb51000011010,adb51000011011,adb51000011100,adb51000011101,adb51000011110,adb51000011111,adb51000100000,adb51000100001,adb51000100010,adb51000100011,adb51000100100,adb51000100101,adb51000100110,adb51000100111,adb51000101000,adb51000101001,adb51000101010,adb51000101011,adb51000101100,adb51000101101,adb51000101110,adb51000101111,adb51000110000,adb51000110001,adb51000110010,adb51000110011,adb51000110100,adb51000110101,adb51000110110,adb51000110111,adb51000111000,adb51000111001,adb51000111010,adb51000111011,adb51000111100,adb51000111101,adb51000111110,adb51000111111,adb51001000000,adb51001000001,adb51001000010,adb51001000011,adb51001000100,adb51001000101,adb51001000110,adb51001000111,adb51001001000,adb51001001001,adb51001001010,adb51001001011,adb51001001100,adb51001001101,adb51001001110,adb51001001111,adb51001010000,adb51001010001,adb51001010010,adb51001010011,adb51001010100,adb51001010101,adb51001010110,adb51001010111,adb51001011000,adb51001011001,adb51001011010,adb51001011011,adb51001011100,adb51001011101,adb51001011110,adb51001011111,adb51001100000,adb51001100001,adb51001100010,adb51001100011,adb51001100100,adb51001100101,adb51001100110,adb51001100111,adb51001101000,adb51001101001,adb51001101010,adb51001101011,adb51001101100,adb51001101101,adb51001101110,adb51001101111,adb51001110000,adb51001110001,adb51001110010,adb51001110011,adb51001110100,adb51001110101,adb51001110110,adb51001110111,adb51001111000,adb51001111001,adb51001111010,adb51001111011,adb51001111100,adb51001111101,adb51001111110,adb51001111111,adb51010000000,adb51010000001,adb51010000010,adb51010000011,adb51010000100,adb51010000101,adb51010000110,adb51010000111,adb51010001000,adb51010001001,adb51010001010,adb51010001011,adb51010001100,adb51010001101,adb51010001110,adb51010001111,adb51010010000,adb51010010001,adb51010010010,adb51010010011,adb51010010100,adb51010010101,adb51010010110,adb51010010111,adb51010011000,adb51010011001,adb51010011010,adb51010011011,adb51010011100,adb51010011101,adb51010011110,adb51010011111,adb51010100000,adb51010100001,adb51010100010,adb51010100011,adb51010100100,adb51010100101,adb51010100110,adb51010100111,adb51010101000,adb51010101001,adb51010101010,adb51010101011,adb51010101100,adb51010101101,adb51010101110,adb51010101111,adb51010110000,adb51010110001,adb51010110010,adb51010110011,adb51010110100,adb51010110101,adb51010110110,adb51010110111,adb51010111000,adb51010111001,adb51010111010,adb51010111011,adb51010111100,adb51010111101,adb51010111110,adb51010111111,adb51011000000,adb51011000001,adb51011000010,adb51011000011,adb51011000100,adb51011000101,adb51011000110,adb51011000111,adb51011001000,adb51011001001,adb51011001010,adb51011001011,adb51011001100,adb51011001101,adb51011001110,adb51011001111,adb51011010000,adb51011010001,adb51011010010,adb51011010011,adb51011010100,adb51011010101,adb51011010110,adb51011010111,adb51011011000,adb51011011001,adb51011011010,adb51011011011,adb51011011100,adb51011011101,adb51011011110,adb51011011111,adb51011100000,adb51011100001,adb51011100010,adb51011100011,adb51011100100,adb51011100101,adb51011100110,adb51011100111,adb51011101000,adb51011101001,adb51011101010,adb51011101011,adb51011101100,adb51011101101,adb51011101110,adb51011101111,adb51011110000,adb51011110001,adb51011110010,adb51011110011,adb51011110100,adb51011110101,adb51011110110,adb51011110111,adb51011111000,adb51011111001,adb51011111010,adb51011111011,adb51011111100,adb51011111101,adb51011111110,adb51011111111,adb51100000000,adb51100000001,adb51100000010,adb51100000011,adb51100000100,adb51100000101,adb51100000110,adb51100000111,adb51100001000,adb51100001001,adb51100001010,adb51100001011,adb51100001100,adb51100001101,adb51100001110,adb51100001111,adb51100010000,adb51100010001,adb51100010010,adb51100010011,adb51100010100,adb51100010101,adb51100010110,adb51100010111,adb51100011000,adb51100011001,adb51100011010,adb51100011011,adb51100011100,adb51100011101,adb51100011110,adb51100011111,adb51100100000,adb51100100001,adb51100100010,adb51100100011,adb51100100100,adb51100100101,adb51100100110,adb51100100111,adb51100101000,adb51100101001,adb51100101010,adb51100101011,adb51100101100,adb51100101101,adb51100101110,adb51100101111,adb51100110000,adb51100110001,adb51100110010,adb51100110011,adb51100110100,adb51100110101,adb51100110110,adb51100110111,adb51100111000,adb51100111001,adb51100111010,adb51100111011,adb51100111100,adb51100111101,adb51100111110,adb51100111111,adb51101000000,adb51101000001,adb51101000010,adb51101000011,adb51101000100,adb51101000101,adb51101000110,adb51101000111,adb51101001000,adb51101001001,adb51101001010,adb51101001011,adb51101001100,adb51101001101,adb51101001110,adb51101001111,adb51101010000,adb51101010001,adb51101010010,adb51101010011,adb51101010100,adb51101010101,adb51101010110,adb51101010111,adb51101011000,adb51101011001,adb51101011010,adb51101011011,adb51101011100,adb51101011101,adb51101011110,adb51101011111,adb51101100000,adb51101100001,adb51101100010,adb51101100011,adb51101100100,adb51101100101,adb51101100110,adb51101100111,adb51101101000,adb51101101001,adb51101101010,adb51101101011,adb51101101100,adb51101101101,adb51101101110,adb51101101111,adb51101110000,adb51101110001,adb51101110010,adb51101110011,adb51101110100,adb51101110101,adb51101110110,adb51101110111,adb51101111000,adb51101111001,adb51101111010,adb51101111011,adb51101111100,adb51101111101,adb51101111110,adb51101111111,adb51110000000,adb51110000001,adb51110000010,adb51110000011,adb51110000100,adb51110000101,adb51110000110,adb51110000111,adb51110001000,adb51110001001,adb51110001010,adb51110001011,adb51110001100,adb51110001101,adb51110001110,adb51110001111,adb51110010000,adb51110010001,adb51110010010,adb51110010011,adb51110010100,adb51110010101,adb51110010110,adb51110010111,adb51110011000,adb51110011001,adb51110011010,adb51110011011,adb51110011100,adb51110011101,adb51110011110,adb51110011111,adb51110100000,adb51110100001,adb51110100010,adb51110100011,adb51110100100,adb51110100101,adb51110100110,adb51110100111,adb51110101000,adb51110101001,adb51110101010,adb51110101011,adb51110101100,adb51110101101,adb51110101110,adb51110101111,adb51110110000,adb51110110001,adb51110110010,adb51110110011,adb51110110100,adb51110110101,adb51110110110,adb51110110111,adb51110111000,adb51110111001,adb51110111010,adb51110111011,adb51110111100,adb51110111101,adb51110111110,adb51110111111,adb51111000000,adb51111000001,adb51111000010,adb51111000011,adb51111000100,adb51111000101,adb51111000110,adb51111000111,adb51111001000,adb51111001001,adb51111001010,adb51111001011,adb51111001100,adb51111001101,adb51111001110,adb51111001111,adb51111010000,adb51111010001,adb51111010010,adb51111010011,adb51111010100,adb51111010101,adb51111010110,adb51111010111,adb51111011000,adb51111011001,adb51111011010,adb51111011011,adb51111011100,adb51111011101,adb51111011110,adb51111011111,adb51111100000,adb51111100001,adb51111100010,adb51111100011,adb51111100100,adb51111100101,adb51111100110,adb51111100111,adb51111101000,adb51111101001,adb51111101010,adb51111101011,adb51111101100,adb51111101101,adb51111101110,adb51111101111,adb51111110000,adb51111110001,adb51111110010,adb51111110011,adb51111110100,adb51111110101,adb51111110110,adb51111110111,adb51111111000,adb51111111001,adb51111111010,adb51111111011,adb51111111100,adb51111111101,adb51111111110,adb51111111111,adbp102,adbp110,adbp118,adbp126,adbp134,adbp142,adbp150,adbp158,adbp202,adbp210,adbp218,adbp226,adbp234,adbp242,adbp250,adbp258),
       Db6(db6,adb600,adb601,adb610,adb611,adb60000000000,adb60000000001,adb60000000010,adb60000000011,adb60000000100,adb60000000101,adb60000000110,adb60000000111,adb60000001000,adb60000001001,adb60000001010,adb60000001011,adb60000001100,adb60000001101,adb60000001110,adb60000001111,adb60000010000,adb60000010001,adb60000010010,adb60000010011,adb60000010100,adb60000010101,adb60000010110,adb60000010111,adb60000011000,adb60000011001,adb60000011010,adb60000011011,adb60000011100,adb60000011101,adb60000011110,adb60000011111,adb60000100000,adb60000100001,adb60000100010,adb60000100011,adb60000100100,adb60000100101,adb60000100110,adb60000100111,adb60000101000,adb60000101001,adb60000101010,adb60000101011,adb60000101100,adb60000101101,adb60000101110,adb60000101111,adb60000110000,adb60000110001,adb60000110010,adb60000110011,adb60000110100,adb60000110101,adb60000110110,adb60000110111,adb60000111000,adb60000111001,adb60000111010,adb60000111011,adb60000111100,adb60000111101,adb60000111110,adb60000111111,adb60001000000,adb60001000001,adb60001000010,adb60001000011,adb60001000100,adb60001000101,adb60001000110,adb60001000111,adb60001001000,adb60001001001,adb60001001010,adb60001001011,adb60001001100,adb60001001101,adb60001001110,adb60001001111,adb60001010000,adb60001010001,adb60001010010,adb60001010011,adb60001010100,adb60001010101,adb60001010110,adb60001010111,adb60001011000,adb60001011001,adb60001011010,adb60001011011,adb60001011100,adb60001011101,adb60001011110,adb60001011111,adb60001100000,adb60001100001,adb60001100010,adb60001100011,adb60001100100,adb60001100101,adb60001100110,adb60001100111,adb60001101000,adb60001101001,adb60001101010,adb60001101011,adb60001101100,adb60001101101,adb60001101110,adb60001101111,adb60001110000,adb60001110001,adb60001110010,adb60001110011,adb60001110100,adb60001110101,adb60001110110,adb60001110111,adb60001111000,adb60001111001,adb60001111010,adb60001111011,adb60001111100,adb60001111101,adb60001111110,adb60001111111,adb60010000000,adb60010000001,adb60010000010,adb60010000011,adb60010000100,adb60010000101,adb60010000110,adb60010000111,adb60010001000,adb60010001001,adb60010001010,adb60010001011,adb60010001100,adb60010001101,adb60010001110,adb60010001111,adb60010010000,adb60010010001,adb60010010010,adb60010010011,adb60010010100,adb60010010101,adb60010010110,adb60010010111,adb60010011000,adb60010011001,adb60010011010,adb60010011011,adb60010011100,adb60010011101,adb60010011110,adb60010011111,adb60010100000,adb60010100001,adb60010100010,adb60010100011,adb60010100100,adb60010100101,adb60010100110,adb60010100111,adb60010101000,adb60010101001,adb60010101010,adb60010101011,adb60010101100,adb60010101101,adb60010101110,adb60010101111,adb60010110000,adb60010110001,adb60010110010,adb60010110011,adb60010110100,adb60010110101,adb60010110110,adb60010110111,adb60010111000,adb60010111001,adb60010111010,adb60010111011,adb60010111100,adb60010111101,adb60010111110,adb60010111111,adb60011000000,adb60011000001,adb60011000010,adb60011000011,adb60011000100,adb60011000101,adb60011000110,adb60011000111,adb60011001000,adb60011001001,adb60011001010,adb60011001011,adb60011001100,adb60011001101,adb60011001110,adb60011001111,adb60011010000,adb60011010001,adb60011010010,adb60011010011,adb60011010100,adb60011010101,adb60011010110,adb60011010111,adb60011011000,adb60011011001,adb60011011010,adb60011011011,adb60011011100,adb60011011101,adb60011011110,adb60011011111,adb60011100000,adb60011100001,adb60011100010,adb60011100011,adb60011100100,adb60011100101,adb60011100110,adb60011100111,adb60011101000,adb60011101001,adb60011101010,adb60011101011,adb60011101100,adb60011101101,adb60011101110,adb60011101111,adb60011110000,adb60011110001,adb60011110010,adb60011110011,adb60011110100,adb60011110101,adb60011110110,adb60011110111,adb60011111000,adb60011111001,adb60011111010,adb60011111011,adb60011111100,adb60011111101,adb60011111110,adb60011111111,adb60100000000,adb60100000001,adb60100000010,adb60100000011,adb60100000100,adb60100000101,adb60100000110,adb60100000111,adb60100001000,adb60100001001,adb60100001010,adb60100001011,adb60100001100,adb60100001101,adb60100001110,adb60100001111,adb60100010000,adb60100010001,adb60100010010,adb60100010011,adb60100010100,adb60100010101,adb60100010110,adb60100010111,adb60100011000,adb60100011001,adb60100011010,adb60100011011,adb60100011100,adb60100011101,adb60100011110,adb60100011111,adb60100100000,adb60100100001,adb60100100010,adb60100100011,adb60100100100,adb60100100101,adb60100100110,adb60100100111,adb60100101000,adb60100101001,adb60100101010,adb60100101011,adb60100101100,adb60100101101,adb60100101110,adb60100101111,adb60100110000,adb60100110001,adb60100110010,adb60100110011,adb60100110100,adb60100110101,adb60100110110,adb60100110111,adb60100111000,adb60100111001,adb60100111010,adb60100111011,adb60100111100,adb60100111101,adb60100111110,adb60100111111,adb60101000000,adb60101000001,adb60101000010,adb60101000011,adb60101000100,adb60101000101,adb60101000110,adb60101000111,adb60101001000,adb60101001001,adb60101001010,adb60101001011,adb60101001100,adb60101001101,adb60101001110,adb60101001111,adb60101010000,adb60101010001,adb60101010010,adb60101010011,adb60101010100,adb60101010101,adb60101010110,adb60101010111,adb60101011000,adb60101011001,adb60101011010,adb60101011011,adb60101011100,adb60101011101,adb60101011110,adb60101011111,adb60101100000,adb60101100001,adb60101100010,adb60101100011,adb60101100100,adb60101100101,adb60101100110,adb60101100111,adb60101101000,adb60101101001,adb60101101010,adb60101101011,adb60101101100,adb60101101101,adb60101101110,adb60101101111,adb60101110000,adb60101110001,adb60101110010,adb60101110011,adb60101110100,adb60101110101,adb60101110110,adb60101110111,adb60101111000,adb60101111001,adb60101111010,adb60101111011,adb60101111100,adb60101111101,adb60101111110,adb60101111111,adb60110000000,adb60110000001,adb60110000010,adb60110000011,adb60110000100,adb60110000101,adb60110000110,adb60110000111,adb60110001000,adb60110001001,adb60110001010,adb60110001011,adb60110001100,adb60110001101,adb60110001110,adb60110001111,adb60110010000,adb60110010001,adb60110010010,adb60110010011,adb60110010100,adb60110010101,adb60110010110,adb60110010111,adb60110011000,adb60110011001,adb60110011010,adb60110011011,adb60110011100,adb60110011101,adb60110011110,adb60110011111,adb60110100000,adb60110100001,adb60110100010,adb60110100011,adb60110100100,adb60110100101,adb60110100110,adb60110100111,adb60110101000,adb60110101001,adb60110101010,adb60110101011,adb60110101100,adb60110101101,adb60110101110,adb60110101111,adb60110110000,adb60110110001,adb60110110010,adb60110110011,adb60110110100,adb60110110101,adb60110110110,adb60110110111,adb60110111000,adb60110111001,adb60110111010,adb60110111011,adb60110111100,adb60110111101,adb60110111110,adb60110111111,adb60111000000,adb60111000001,adb60111000010,adb60111000011,adb60111000100,adb60111000101,adb60111000110,adb60111000111,adb60111001000,adb60111001001,adb60111001010,adb60111001011,adb60111001100,adb60111001101,adb60111001110,adb60111001111,adb60111010000,adb60111010001,adb60111010010,adb60111010011,adb60111010100,adb60111010101,adb60111010110,adb60111010111,adb60111011000,adb60111011001,adb60111011010,adb60111011011,adb60111011100,adb60111011101,adb60111011110,adb60111011111,adb60111100000,adb60111100001,adb60111100010,adb60111100011,adb60111100100,adb60111100101,adb60111100110,adb60111100111,adb60111101000,adb60111101001,adb60111101010,adb60111101011,adb60111101100,adb60111101101,adb60111101110,adb60111101111,adb60111110000,adb60111110001,adb60111110010,adb60111110011,adb60111110100,adb60111110101,adb60111110110,adb60111110111,adb60111111000,adb60111111001,adb60111111010,adb60111111011,adb60111111100,adb60111111101,adb60111111110,adb60111111111,adb61000000000,adb61000000001,adb61000000010,adb61000000011,adb61000000100,adb61000000101,adb61000000110,adb61000000111,adb61000001000,adb61000001001,adb61000001010,adb61000001011,adb61000001100,adb61000001101,adb61000001110,adb61000001111,adb61000010000,adb61000010001,adb61000010010,adb61000010011,adb61000010100,adb61000010101,adb61000010110,adb61000010111,adb61000011000,adb61000011001,adb61000011010,adb61000011011,adb61000011100,adb61000011101,adb61000011110,adb61000011111,adb61000100000,adb61000100001,adb61000100010,adb61000100011,adb61000100100,adb61000100101,adb61000100110,adb61000100111,adb61000101000,adb61000101001,adb61000101010,adb61000101011,adb61000101100,adb61000101101,adb61000101110,adb61000101111,adb61000110000,adb61000110001,adb61000110010,adb61000110011,adb61000110100,adb61000110101,adb61000110110,adb61000110111,adb61000111000,adb61000111001,adb61000111010,adb61000111011,adb61000111100,adb61000111101,adb61000111110,adb61000111111,adb61001000000,adb61001000001,adb61001000010,adb61001000011,adb61001000100,adb61001000101,adb61001000110,adb61001000111,adb61001001000,adb61001001001,adb61001001010,adb61001001011,adb61001001100,adb61001001101,adb61001001110,adb61001001111,adb61001010000,adb61001010001,adb61001010010,adb61001010011,adb61001010100,adb61001010101,adb61001010110,adb61001010111,adb61001011000,adb61001011001,adb61001011010,adb61001011011,adb61001011100,adb61001011101,adb61001011110,adb61001011111,adb61001100000,adb61001100001,adb61001100010,adb61001100011,adb61001100100,adb61001100101,adb61001100110,adb61001100111,adb61001101000,adb61001101001,adb61001101010,adb61001101011,adb61001101100,adb61001101101,adb61001101110,adb61001101111,adb61001110000,adb61001110001,adb61001110010,adb61001110011,adb61001110100,adb61001110101,adb61001110110,adb61001110111,adb61001111000,adb61001111001,adb61001111010,adb61001111011,adb61001111100,adb61001111101,adb61001111110,adb61001111111,adb61010000000,adb61010000001,adb61010000010,adb61010000011,adb61010000100,adb61010000101,adb61010000110,adb61010000111,adb61010001000,adb61010001001,adb61010001010,adb61010001011,adb61010001100,adb61010001101,adb61010001110,adb61010001111,adb61010010000,adb61010010001,adb61010010010,adb61010010011,adb61010010100,adb61010010101,adb61010010110,adb61010010111,adb61010011000,adb61010011001,adb61010011010,adb61010011011,adb61010011100,adb61010011101,adb61010011110,adb61010011111,adb61010100000,adb61010100001,adb61010100010,adb61010100011,adb61010100100,adb61010100101,adb61010100110,adb61010100111,adb61010101000,adb61010101001,adb61010101010,adb61010101011,adb61010101100,adb61010101101,adb61010101110,adb61010101111,adb61010110000,adb61010110001,adb61010110010,adb61010110011,adb61010110100,adb61010110101,adb61010110110,adb61010110111,adb61010111000,adb61010111001,adb61010111010,adb61010111011,adb61010111100,adb61010111101,adb61010111110,adb61010111111,adb61011000000,adb61011000001,adb61011000010,adb61011000011,adb61011000100,adb61011000101,adb61011000110,adb61011000111,adb61011001000,adb61011001001,adb61011001010,adb61011001011,adb61011001100,adb61011001101,adb61011001110,adb61011001111,adb61011010000,adb61011010001,adb61011010010,adb61011010011,adb61011010100,adb61011010101,adb61011010110,adb61011010111,adb61011011000,adb61011011001,adb61011011010,adb61011011011,adb61011011100,adb61011011101,adb61011011110,adb61011011111,adb61011100000,adb61011100001,adb61011100010,adb61011100011,adb61011100100,adb61011100101,adb61011100110,adb61011100111,adb61011101000,adb61011101001,adb61011101010,adb61011101011,adb61011101100,adb61011101101,adb61011101110,adb61011101111,adb61011110000,adb61011110001,adb61011110010,adb61011110011,adb61011110100,adb61011110101,adb61011110110,adb61011110111,adb61011111000,adb61011111001,adb61011111010,adb61011111011,adb61011111100,adb61011111101,adb61011111110,adb61011111111,adb61100000000,adb61100000001,adb61100000010,adb61100000011,adb61100000100,adb61100000101,adb61100000110,adb61100000111,adb61100001000,adb61100001001,adb61100001010,adb61100001011,adb61100001100,adb61100001101,adb61100001110,adb61100001111,adb61100010000,adb61100010001,adb61100010010,adb61100010011,adb61100010100,adb61100010101,adb61100010110,adb61100010111,adb61100011000,adb61100011001,adb61100011010,adb61100011011,adb61100011100,adb61100011101,adb61100011110,adb61100011111,adb61100100000,adb61100100001,adb61100100010,adb61100100011,adb61100100100,adb61100100101,adb61100100110,adb61100100111,adb61100101000,adb61100101001,adb61100101010,adb61100101011,adb61100101100,adb61100101101,adb61100101110,adb61100101111,adb61100110000,adb61100110001,adb61100110010,adb61100110011,adb61100110100,adb61100110101,adb61100110110,adb61100110111,adb61100111000,adb61100111001,adb61100111010,adb61100111011,adb61100111100,adb61100111101,adb61100111110,adb61100111111,adb61101000000,adb61101000001,adb61101000010,adb61101000011,adb61101000100,adb61101000101,adb61101000110,adb61101000111,adb61101001000,adb61101001001,adb61101001010,adb61101001011,adb61101001100,adb61101001101,adb61101001110,adb61101001111,adb61101010000,adb61101010001,adb61101010010,adb61101010011,adb61101010100,adb61101010101,adb61101010110,adb61101010111,adb61101011000,adb61101011001,adb61101011010,adb61101011011,adb61101011100,adb61101011101,adb61101011110,adb61101011111,adb61101100000,adb61101100001,adb61101100010,adb61101100011,adb61101100100,adb61101100101,adb61101100110,adb61101100111,adb61101101000,adb61101101001,adb61101101010,adb61101101011,adb61101101100,adb61101101101,adb61101101110,adb61101101111,adb61101110000,adb61101110001,adb61101110010,adb61101110011,adb61101110100,adb61101110101,adb61101110110,adb61101110111,adb61101111000,adb61101111001,adb61101111010,adb61101111011,adb61101111100,adb61101111101,adb61101111110,adb61101111111,adb61110000000,adb61110000001,adb61110000010,adb61110000011,adb61110000100,adb61110000101,adb61110000110,adb61110000111,adb61110001000,adb61110001001,adb61110001010,adb61110001011,adb61110001100,adb61110001101,adb61110001110,adb61110001111,adb61110010000,adb61110010001,adb61110010010,adb61110010011,adb61110010100,adb61110010101,adb61110010110,adb61110010111,adb61110011000,adb61110011001,adb61110011010,adb61110011011,adb61110011100,adb61110011101,adb61110011110,adb61110011111,adb61110100000,adb61110100001,adb61110100010,adb61110100011,adb61110100100,adb61110100101,adb61110100110,adb61110100111,adb61110101000,adb61110101001,adb61110101010,adb61110101011,adb61110101100,adb61110101101,adb61110101110,adb61110101111,adb61110110000,adb61110110001,adb61110110010,adb61110110011,adb61110110100,adb61110110101,adb61110110110,adb61110110111,adb61110111000,adb61110111001,adb61110111010,adb61110111011,adb61110111100,adb61110111101,adb61110111110,adb61110111111,adb61111000000,adb61111000001,adb61111000010,adb61111000011,adb61111000100,adb61111000101,adb61111000110,adb61111000111,adb61111001000,adb61111001001,adb61111001010,adb61111001011,adb61111001100,adb61111001101,adb61111001110,adb61111001111,adb61111010000,adb61111010001,adb61111010010,adb61111010011,adb61111010100,adb61111010101,adb61111010110,adb61111010111,adb61111011000,adb61111011001,adb61111011010,adb61111011011,adb61111011100,adb61111011101,adb61111011110,adb61111011111,adb61111100000,adb61111100001,adb61111100010,adb61111100011,adb61111100100,adb61111100101,adb61111100110,adb61111100111,adb61111101000,adb61111101001,adb61111101010,adb61111101011,adb61111101100,adb61111101101,adb61111101110,adb61111101111,adb61111110000,adb61111110001,adb61111110010,adb61111110011,adb61111110100,adb61111110101,adb61111110110,adb61111110111,adb61111111000,adb61111111001,adb61111111010,adb61111111011,adb61111111100,adb61111111101,adb61111111110,adb61111111111,adbp109,adbp117,adbp125,adbp133,adbp141,adbp149,adbp157,adbp209,adbp217,adbp225,adbp233,adbp241,adbp249,adbp257,adbtopline1),
       Db7(db7,adb700,adb701,adb710,adb711,adb70000000000,adb70000000001,adb70000000010,adb70000000011,adb70000000100,adb70000000101,adb70000000110,adb70000000111,adb70000001000,adb70000001001,adb70000001010,adb70000001011,adb70000001100,adb70000001101,adb70000001110,adb70000001111,adb70000010000,adb70000010001,adb70000010010,adb70000010011,adb70000010100,adb70000010101,adb70000010110,adb70000010111,adb70000011000,adb70000011001,adb70000011010,adb70000011011,adb70000011100,adb70000011101,adb70000011110,adb70000011111,adb70000100000,adb70000100001,adb70000100010,adb70000100011,adb70000100100,adb70000100101,adb70000100110,adb70000100111,adb70000101000,adb70000101001,adb70000101010,adb70000101011,adb70000101100,adb70000101101,adb70000101110,adb70000101111,adb70000110000,adb70000110001,adb70000110010,adb70000110011,adb70000110100,adb70000110101,adb70000110110,adb70000110111,adb70000111000,adb70000111001,adb70000111010,adb70000111011,adb70000111100,adb70000111101,adb70000111110,adb70000111111,adb70001000000,adb70001000001,adb70001000010,adb70001000011,adb70001000100,adb70001000101,adb70001000110,adb70001000111,adb70001001000,adb70001001001,adb70001001010,adb70001001011,adb70001001100,adb70001001101,adb70001001110,adb70001001111,adb70001010000,adb70001010001,adb70001010010,adb70001010011,adb70001010100,adb70001010101,adb70001010110,adb70001010111,adb70001011000,adb70001011001,adb70001011010,adb70001011011,adb70001011100,adb70001011101,adb70001011110,adb70001011111,adb70001100000,adb70001100001,adb70001100010,adb70001100011,adb70001100100,adb70001100101,adb70001100110,adb70001100111,adb70001101000,adb70001101001,adb70001101010,adb70001101011,adb70001101100,adb70001101101,adb70001101110,adb70001101111,adb70001110000,adb70001110001,adb70001110010,adb70001110011,adb70001110100,adb70001110101,adb70001110110,adb70001110111,adb70001111000,adb70001111001,adb70001111010,adb70001111011,adb70001111100,adb70001111101,adb70001111110,adb70001111111,adb70010000000,adb70010000001,adb70010000010,adb70010000011,adb70010000100,adb70010000101,adb70010000110,adb70010000111,adb70010001000,adb70010001001,adb70010001010,adb70010001011,adb70010001100,adb70010001101,adb70010001110,adb70010001111,adb70010010000,adb70010010001,adb70010010010,adb70010010011,adb70010010100,adb70010010101,adb70010010110,adb70010010111,adb70010011000,adb70010011001,adb70010011010,adb70010011011,adb70010011100,adb70010011101,adb70010011110,adb70010011111,adb70010100000,adb70010100001,adb70010100010,adb70010100011,adb70010100100,adb70010100101,adb70010100110,adb70010100111,adb70010101000,adb70010101001,adb70010101010,adb70010101011,adb70010101100,adb70010101101,adb70010101110,adb70010101111,adb70010110000,adb70010110001,adb70010110010,adb70010110011,adb70010110100,adb70010110101,adb70010110110,adb70010110111,adb70010111000,adb70010111001,adb70010111010,adb70010111011,adb70010111100,adb70010111101,adb70010111110,adb70010111111,adb70011000000,adb70011000001,adb70011000010,adb70011000011,adb70011000100,adb70011000101,adb70011000110,adb70011000111,adb70011001000,adb70011001001,adb70011001010,adb70011001011,adb70011001100,adb70011001101,adb70011001110,adb70011001111,adb70011010000,adb70011010001,adb70011010010,adb70011010011,adb70011010100,adb70011010101,adb70011010110,adb70011010111,adb70011011000,adb70011011001,adb70011011010,adb70011011011,adb70011011100,adb70011011101,adb70011011110,adb70011011111,adb70011100000,adb70011100001,adb70011100010,adb70011100011,adb70011100100,adb70011100101,adb70011100110,adb70011100111,adb70011101000,adb70011101001,adb70011101010,adb70011101011,adb70011101100,adb70011101101,adb70011101110,adb70011101111,adb70011110000,adb70011110001,adb70011110010,adb70011110011,adb70011110100,adb70011110101,adb70011110110,adb70011110111,adb70011111000,adb70011111001,adb70011111010,adb70011111011,adb70011111100,adb70011111101,adb70011111110,adb70011111111,adb70100000000,adb70100000001,adb70100000010,adb70100000011,adb70100000100,adb70100000101,adb70100000110,adb70100000111,adb70100001000,adb70100001001,adb70100001010,adb70100001011,adb70100001100,adb70100001101,adb70100001110,adb70100001111,adb70100010000,adb70100010001,adb70100010010,adb70100010011,adb70100010100,adb70100010101,adb70100010110,adb70100010111,adb70100011000,adb70100011001,adb70100011010,adb70100011011,adb70100011100,adb70100011101,adb70100011110,adb70100011111,adb70100100000,adb70100100001,adb70100100010,adb70100100011,adb70100100100,adb70100100101,adb70100100110,adb70100100111,adb70100101000,adb70100101001,adb70100101010,adb70100101011,adb70100101100,adb70100101101,adb70100101110,adb70100101111,adb70100110000,adb70100110001,adb70100110010,adb70100110011,adb70100110100,adb70100110101,adb70100110110,adb70100110111,adb70100111000,adb70100111001,adb70100111010,adb70100111011,adb70100111100,adb70100111101,adb70100111110,adb70100111111,adb70101000000,adb70101000001,adb70101000010,adb70101000011,adb70101000100,adb70101000101,adb70101000110,adb70101000111,adb70101001000,adb70101001001,adb70101001010,adb70101001011,adb70101001100,adb70101001101,adb70101001110,adb70101001111,adb70101010000,adb70101010001,adb70101010010,adb70101010011,adb70101010100,adb70101010101,adb70101010110,adb70101010111,adb70101011000,adb70101011001,adb70101011010,adb70101011011,adb70101011100,adb70101011101,adb70101011110,adb70101011111,adb70101100000,adb70101100001,adb70101100010,adb70101100011,adb70101100100,adb70101100101,adb70101100110,adb70101100111,adb70101101000,adb70101101001,adb70101101010,adb70101101011,adb70101101100,adb70101101101,adb70101101110,adb70101101111,adb70101110000,adb70101110001,adb70101110010,adb70101110011,adb70101110100,adb70101110101,adb70101110110,adb70101110111,adb70101111000,adb70101111001,adb70101111010,adb70101111011,adb70101111100,adb70101111101,adb70101111110,adb70101111111,adb70110000000,adb70110000001,adb70110000010,adb70110000011,adb70110000100,adb70110000101,adb70110000110,adb70110000111,adb70110001000,adb70110001001,adb70110001010,adb70110001011,adb70110001100,adb70110001101,adb70110001110,adb70110001111,adb70110010000,adb70110010001,adb70110010010,adb70110010011,adb70110010100,adb70110010101,adb70110010110,adb70110010111,adb70110011000,adb70110011001,adb70110011010,adb70110011011,adb70110011100,adb70110011101,adb70110011110,adb70110011111,adb70110100000,adb70110100001,adb70110100010,adb70110100011,adb70110100100,adb70110100101,adb70110100110,adb70110100111,adb70110101000,adb70110101001,adb70110101010,adb70110101011,adb70110101100,adb70110101101,adb70110101110,adb70110101111,adb70110110000,adb70110110001,adb70110110010,adb70110110011,adb70110110100,adb70110110101,adb70110110110,adb70110110111,adb70110111000,adb70110111001,adb70110111010,adb70110111011,adb70110111100,adb70110111101,adb70110111110,adb70110111111,adb70111000000,adb70111000001,adb70111000010,adb70111000011,adb70111000100,adb70111000101,adb70111000110,adb70111000111,adb70111001000,adb70111001001,adb70111001010,adb70111001011,adb70111001100,adb70111001101,adb70111001110,adb70111001111,adb70111010000,adb70111010001,adb70111010010,adb70111010011,adb70111010100,adb70111010101,adb70111010110,adb70111010111,adb70111011000,adb70111011001,adb70111011010,adb70111011011,adb70111011100,adb70111011101,adb70111011110,adb70111011111,adb70111100000,adb70111100001,adb70111100010,adb70111100011,adb70111100100,adb70111100101,adb70111100110,adb70111100111,adb70111101000,adb70111101001,adb70111101010,adb70111101011,adb70111101100,adb70111101101,adb70111101110,adb70111101111,adb70111110000,adb70111110001,adb70111110010,adb70111110011,adb70111110100,adb70111110101,adb70111110110,adb70111110111,adb70111111000,adb70111111001,adb70111111010,adb70111111011,adb70111111100,adb70111111101,adb70111111110,adb70111111111,adb71000000000,adb71000000001,adb71000000010,adb71000000011,adb71000000100,adb71000000101,adb71000000110,adb71000000111,adb71000001000,adb71000001001,adb71000001010,adb71000001011,adb71000001100,adb71000001101,adb71000001110,adb71000001111,adb71000010000,adb71000010001,adb71000010010,adb71000010011,adb71000010100,adb71000010101,adb71000010110,adb71000010111,adb71000011000,adb71000011001,adb71000011010,adb71000011011,adb71000011100,adb71000011101,adb71000011110,adb71000011111,adb71000100000,adb71000100001,adb71000100010,adb71000100011,adb71000100100,adb71000100101,adb71000100110,adb71000100111,adb71000101000,adb71000101001,adb71000101010,adb71000101011,adb71000101100,adb71000101101,adb71000101110,adb71000101111,adb71000110000,adb71000110001,adb71000110010,adb71000110011,adb71000110100,adb71000110101,adb71000110110,adb71000110111,adb71000111000,adb71000111001,adb71000111010,adb71000111011,adb71000111100,adb71000111101,adb71000111110,adb71000111111,adb71001000000,adb71001000001,adb71001000010,adb71001000011,adb71001000100,adb71001000101,adb71001000110,adb71001000111,adb71001001000,adb71001001001,adb71001001010,adb71001001011,adb71001001100,adb71001001101,adb71001001110,adb71001001111,adb71001010000,adb71001010001,adb71001010010,adb71001010011,adb71001010100,adb71001010101,adb71001010110,adb71001010111,adb71001011000,adb71001011001,adb71001011010,adb71001011011,adb71001011100,adb71001011101,adb71001011110,adb71001011111,adb71001100000,adb71001100001,adb71001100010,adb71001100011,adb71001100100,adb71001100101,adb71001100110,adb71001100111,adb71001101000,adb71001101001,adb71001101010,adb71001101011,adb71001101100,adb71001101101,adb71001101110,adb71001101111,adb71001110000,adb71001110001,adb71001110010,adb71001110011,adb71001110100,adb71001110101,adb71001110110,adb71001110111,adb71001111000,adb71001111001,adb71001111010,adb71001111011,adb71001111100,adb71001111101,adb71001111110,adb71001111111,adb71010000000,adb71010000001,adb71010000010,adb71010000011,adb71010000100,adb71010000101,adb71010000110,adb71010000111,adb71010001000,adb71010001001,adb71010001010,adb71010001011,adb71010001100,adb71010001101,adb71010001110,adb71010001111,adb71010010000,adb71010010001,adb71010010010,adb71010010011,adb71010010100,adb71010010101,adb71010010110,adb71010010111,adb71010011000,adb71010011001,adb71010011010,adb71010011011,adb71010011100,adb71010011101,adb71010011110,adb71010011111,adb71010100000,adb71010100001,adb71010100010,adb71010100011,adb71010100100,adb71010100101,adb71010100110,adb71010100111,adb71010101000,adb71010101001,adb71010101010,adb71010101011,adb71010101100,adb71010101101,adb71010101110,adb71010101111,adb71010110000,adb71010110001,adb71010110010,adb71010110011,adb71010110100,adb71010110101,adb71010110110,adb71010110111,adb71010111000,adb71010111001,adb71010111010,adb71010111011,adb71010111100,adb71010111101,adb71010111110,adb71010111111,adb71011000000,adb71011000001,adb71011000010,adb71011000011,adb71011000100,adb71011000101,adb71011000110,adb71011000111,adb71011001000,adb71011001001,adb71011001010,adb71011001011,adb71011001100,adb71011001101,adb71011001110,adb71011001111,adb71011010000,adb71011010001,adb71011010010,adb71011010011,adb71011010100,adb71011010101,adb71011010110,adb71011010111,adb71011011000,adb71011011001,adb71011011010,adb71011011011,adb71011011100,adb71011011101,adb71011011110,adb71011011111,adb71011100000,adb71011100001,adb71011100010,adb71011100011,adb71011100100,adb71011100101,adb71011100110,adb71011100111,adb71011101000,adb71011101001,adb71011101010,adb71011101011,adb71011101100,adb71011101101,adb71011101110,adb71011101111,adb71011110000,adb71011110001,adb71011110010,adb71011110011,adb71011110100,adb71011110101,adb71011110110,adb71011110111,adb71011111000,adb71011111001,adb71011111010,adb71011111011,adb71011111100,adb71011111101,adb71011111110,adb71011111111,adb71100000000,adb71100000001,adb71100000010,adb71100000011,adb71100000100,adb71100000101,adb71100000110,adb71100000111,adb71100001000,adb71100001001,adb71100001010,adb71100001011,adb71100001100,adb71100001101,adb71100001110,adb71100001111,adb71100010000,adb71100010001,adb71100010010,adb71100010011,adb71100010100,adb71100010101,adb71100010110,adb71100010111,adb71100011000,adb71100011001,adb71100011010,adb71100011011,adb71100011100,adb71100011101,adb71100011110,adb71100011111,adb71100100000,adb71100100001,adb71100100010,adb71100100011,adb71100100100,adb71100100101,adb71100100110,adb71100100111,adb71100101000,adb71100101001,adb71100101010,adb71100101011,adb71100101100,adb71100101101,adb71100101110,adb71100101111,adb71100110000,adb71100110001,adb71100110010,adb71100110011,adb71100110100,adb71100110101,adb71100110110,adb71100110111,adb71100111000,adb71100111001,adb71100111010,adb71100111011,adb71100111100,adb71100111101,adb71100111110,adb71100111111,adb71101000000,adb71101000001,adb71101000010,adb71101000011,adb71101000100,adb71101000101,adb71101000110,adb71101000111,adb71101001000,adb71101001001,adb71101001010,adb71101001011,adb71101001100,adb71101001101,adb71101001110,adb71101001111,adb71101010000,adb71101010001,adb71101010010,adb71101010011,adb71101010100,adb71101010101,adb71101010110,adb71101010111,adb71101011000,adb71101011001,adb71101011010,adb71101011011,adb71101011100,adb71101011101,adb71101011110,adb71101011111,adb71101100000,adb71101100001,adb71101100010,adb71101100011,adb71101100100,adb71101100101,adb71101100110,adb71101100111,adb71101101000,adb71101101001,adb71101101010,adb71101101011,adb71101101100,adb71101101101,adb71101101110,adb71101101111,adb71101110000,adb71101110001,adb71101110010,adb71101110011,adb71101110100,adb71101110101,adb71101110110,adb71101110111,adb71101111000,adb71101111001,adb71101111010,adb71101111011,adb71101111100,adb71101111101,adb71101111110,adb71101111111,adb71110000000,adb71110000001,adb71110000010,adb71110000011,adb71110000100,adb71110000101,adb71110000110,adb71110000111,adb71110001000,adb71110001001,adb71110001010,adb71110001011,adb71110001100,adb71110001101,adb71110001110,adb71110001111,adb71110010000,adb71110010001,adb71110010010,adb71110010011,adb71110010100,adb71110010101,adb71110010110,adb71110010111,adb71110011000,adb71110011001,adb71110011010,adb71110011011,adb71110011100,adb71110011101,adb71110011110,adb71110011111,adb71110100000,adb71110100001,adb71110100010,adb71110100011,adb71110100100,adb71110100101,adb71110100110,adb71110100111,adb71110101000,adb71110101001,adb71110101010,adb71110101011,adb71110101100,adb71110101101,adb71110101110,adb71110101111,adb71110110000,adb71110110001,adb71110110010,adb71110110011,adb71110110100,adb71110110101,adb71110110110,adb71110110111,adb71110111000,adb71110111001,adb71110111010,adb71110111011,adb71110111100,adb71110111101,adb71110111110,adb71110111111,adb71111000000,adb71111000001,adb71111000010,adb71111000011,adb71111000100,adb71111000101,adb71111000110,adb71111000111,adb71111001000,adb71111001001,adb71111001010,adb71111001011,adb71111001100,adb71111001101,adb71111001110,adb71111001111,adb71111010000,adb71111010001,adb71111010010,adb71111010011,adb71111010100,adb71111010101,adb71111010110,adb71111010111,adb71111011000,adb71111011001,adb71111011010,adb71111011011,adb71111011100,adb71111011101,adb71111011110,adb71111011111,adb71111100000,adb71111100001,adb71111100010,adb71111100011,adb71111100100,adb71111100101,adb71111100110,adb71111100111,adb71111101000,adb71111101001,adb71111101010,adb71111101011,adb71111101100,adb71111101101,adb71111101110,adb71111101111,adb71111110000,adb71111110001,adb71111110010,adb71111110011,adb71111110100,adb71111110101,adb71111110110,adb71111110111,adb71111111000,adb71111111001,adb71111111010,adb71111111011,adb71111111100,adb71111111101,adb71111111110,adb71111111111,adbp108,adbp116,adbp124,adbp132,adbp140,adbp148,adbp156,adbp208,adbp216,adbp224,adbp232,adbp240,adbp248,adbp256,adbtopline1);

and    Adb000(adb000,n0011,n0010,n0009,dbv1),
       Adb001(adb001,n0011,n0010,m0009,dbv0),
       Adb010(adb010,n0011,m0010,n0009,m0017),
       Adb011(adb011,n0011,m0010,m0009,dbv0),
Adb00000000000	(	adb00000000000,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m111111_0	),
Adb00000000001	(	adb00000000001,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m111111_0	),
Adb00000000010	(	adb00000000010,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m111111_0	),
Adb00000000011	(	adb00000000011,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m111111_0	),
Adb00000000100	(	adb00000000100,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m111111_0	),
Adb00000000101	(	adb00000000101,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m111111_0	),
Adb00000000110	(	adb00000000110,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m111111_0	),
Adb00000000111	(	adb00000000111,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m111111_0	),
Adb00000001000	(	adb00000001000,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m111111_0	),
Adb00000001001	(	adb00000001001,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m111111_0	),
Adb00000001010	(	adb00000001010,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m111111_0	),
Adb00000001011	(	adb00000001011,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m111111_0	),
Adb00000001100	(	adb00000001100,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m111111_0	),
Adb00000001101	(	adb00000001101,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m111111_0	),
Adb00000001110	(	adb00000001110,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m111111_0	),
Adb00000001111	(	adb00000001111,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m111111_0	),
Adb00000010000	(	adb00000010000,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m111111_0	),
Adb00000010001	(	adb00000010001,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m111111_0	),
Adb00000010010	(	adb00000010010,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m111111_0	),
Adb00000010011	(	adb00000010011,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m111111_0	),
Adb00000010100	(	adb00000010100,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m111111_0	),
Adb00000010101	(	adb00000010101,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m111111_0	),
Adb00000010110	(	adb00000010110,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m111111_0	),
Adb00000010111	(	adb00000010111,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m111111_0	),
Adb00000011000	(	adb00000011000,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m111111_0	),
Adb00000011001	(	adb00000011001,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m111111_0	),
Adb00000011010	(	adb00000011010,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m111111_0	),
Adb00000011011	(	adb00000011011,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m111111_0	),
Adb00000011100	(	adb00000011100,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m111111_0	),
Adb00000011101	(	adb00000011101,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m111111_0	),
Adb00000011110	(	adb00000011110,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m111111_0	),
Adb00000011111	(	adb00000011111,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m111111_0	),
Adb00000100000	(	adb00000100000,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m111111_0	),
Adb00000100001	(	adb00000100001,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m111111_0	),
Adb00000100010	(	adb00000100010,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m111111_0	),
Adb00000100011	(	adb00000100011,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m111111_0	),
Adb00000100100	(	adb00000100100,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m111111_0	),
Adb00000100101	(	adb00000100101,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m111111_0	),
Adb00000100110	(	adb00000100110,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m111111_0	),
Adb00000100111	(	adb00000100111,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m111111_0	),
Adb00000101000	(	adb00000101000,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m111111_0	),
Adb00000101001	(	adb00000101001,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m111111_0	),
Adb00000101010	(	adb00000101010,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m111111_0	),
Adb00000101011	(	adb00000101011,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m111111_0	),
Adb00000101100	(	adb00000101100,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m111111_0	),
Adb00000101101	(	adb00000101101,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m111111_0	),
Adb00000101110	(	adb00000101110,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m111111_0	),
Adb00000101111	(	adb00000101111,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m111111_0	),
Adb00000110000	(	adb00000110000,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m111111_0	),
Adb00000110001	(	adb00000110001,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m111111_0	),
Adb00000110010	(	adb00000110010,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m111111_0	),
Adb00000110011	(	adb00000110011,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m111111_0	),
Adb00000110100	(	adb00000110100,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m111111_0	),
Adb00000110101	(	adb00000110101,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m111111_0	),
Adb00000110110	(	adb00000110110,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m111111_0	),
Adb00000110111	(	adb00000110111,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m111111_0	),
Adb00000111000	(	adb00000111000,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m111111_0	),
Adb00000111001	(	adb00000111001,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m111111_0	),
Adb00000111010	(	adb00000111010,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m111111_0	),
Adb00000111011	(	adb00000111011,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m111111_0	),
Adb00000111100	(	adb00000111100,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m111111_0	),
Adb00000111101	(	adb00000111101,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m111111_0	),
Adb00000111110	(	adb00000111110,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m111111_0	),
Adb00000111111	(	adb00000111111,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m111111_0	),
Adb00001000000	(	adb00001000000,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m111111_0	),
Adb00001000001	(	adb00001000001,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m111111_0	),
Adb00001000010	(	adb00001000010,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m111111_0	),
Adb00001000011	(	adb00001000011,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m111111_0	),
Adb00001000100	(	adb00001000100,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m111111_0	),
Adb00001000101	(	adb00001000101,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m111111_0	),
Adb00001000110	(	adb00001000110,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m111111_0	),
Adb00001000111	(	adb00001000111,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m111111_0	),
Adb00001001000	(	adb00001001000,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m111111_0	),
Adb00001001001	(	adb00001001001,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m111111_0	),
Adb00001001010	(	adb00001001010,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m111111_0	),
Adb00001001011	(	adb00001001011,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m111111_0	),
Adb00001001100	(	adb00001001100,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m111111_0	),
Adb00001001101	(	adb00001001101,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m111111_0	),
Adb00001001110	(	adb00001001110,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m111111_0	),
Adb00001001111	(	adb00001001111,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m111111_0	),
Adb00001010000	(	adb00001010000,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m111111_0	),
Adb00001010001	(	adb00001010001,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m111111_0	),
Adb00001010010	(	adb00001010010,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m111111_0	),
Adb00001010011	(	adb00001010011,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m111111_0	),
Adb00001010100	(	adb00001010100,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m111111_0	),
Adb00001010101	(	adb00001010101,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m111111_0	),
Adb00001010110	(	adb00001010110,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m111111_0	),
Adb00001010111	(	adb00001010111,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m111111_0	),
Adb00001011000	(	adb00001011000,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m111111_0	),
Adb00001011001	(	adb00001011001,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m111111_0	),
Adb00001011010	(	adb00001011010,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m111111_0	),
Adb00001011011	(	adb00001011011,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m111111_0	),
Adb00001011100	(	adb00001011100,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m111111_0	),
Adb00001011101	(	adb00001011101,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m111111_0	),
Adb00001011110	(	adb00001011110,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m111111_0	),
Adb00001011111	(	adb00001011111,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m111111_0	),
Adb00001100000	(	adb00001100000,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m111111_0	),
Adb00001100001	(	adb00001100001,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m111111_0	),
Adb00001100010	(	adb00001100010,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m111111_0	),
Adb00001100011	(	adb00001100011,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m111111_0	),
Adb00001100100	(	adb00001100100,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m111111_0	),
Adb00001100101	(	adb00001100101,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m111111_0	),
Adb00001100110	(	adb00001100110,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m111111_0	),
Adb00001100111	(	adb00001100111,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m111111_0	),
Adb00001101000	(	adb00001101000,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m111111_0	),
Adb00001101001	(	adb00001101001,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m111111_0	),
Adb00001101010	(	adb00001101010,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m111111_0	),
Adb00001101011	(	adb00001101011,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m111111_0	),
Adb00001101100	(	adb00001101100,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m111111_0	),
Adb00001101101	(	adb00001101101,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m111111_0	),
Adb00001101110	(	adb00001101110,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m111111_0	),
Adb00001101111	(	adb00001101111,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m111111_0	),
Adb00001110000	(	adb00001110000,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m111111_0	),
Adb00001110001	(	adb00001110001,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m111111_0	),
Adb00001110010	(	adb00001110010,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m111111_0	),
Adb00001110011	(	adb00001110011,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m111111_0	),
Adb00001110100	(	adb00001110100,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m111111_0	),
Adb00001110101	(	adb00001110101,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m111111_0	),
Adb00001110110	(	adb00001110110,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m111111_0	),
Adb00001110111	(	adb00001110111,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m111111_0	),
Adb00001111000	(	adb00001111000,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m111111_0	),
Adb00001111001	(	adb00001111001,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m111111_0	),
Adb00001111010	(	adb00001111010,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m111111_0	),
Adb00001111011	(	adb00001111011,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m111111_0	),
Adb00001111100	(	adb00001111100,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m111111_0	),
Adb00001111101	(	adb00001111101,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m111111_0	),
Adb00001111110	(	adb00001111110,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m111111_0	),
Adb00001111111	(	adb00001111111,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m111111_0	),
Adb00010000000	(	adb00010000000,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m110111_0	),
Adb00010000001	(	adb00010000001,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m110111_0	),
Adb00010000010	(	adb00010000010,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m110111_0	),
Adb00010000011	(	adb00010000011,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m110111_0	),
Adb00010000100	(	adb00010000100,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m110111_0	),
Adb00010000101	(	adb00010000101,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m110111_0	),
Adb00010000110	(	adb00010000110,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m110111_0	),
Adb00010000111	(	adb00010000111,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m110111_0	),
Adb00010001000	(	adb00010001000,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m110111_0	),
Adb00010001001	(	adb00010001001,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m110111_0	),
Adb00010001010	(	adb00010001010,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m110111_0	),
Adb00010001011	(	adb00010001011,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m110111_0	),
Adb00010001100	(	adb00010001100,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m110111_0	),
Adb00010001101	(	adb00010001101,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m110111_0	),
Adb00010001110	(	adb00010001110,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m110111_0	),
Adb00010001111	(	adb00010001111,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m110111_0	),
Adb00010010000	(	adb00010010000,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m110111_0	),
Adb00010010001	(	adb00010010001,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m110111_0	),
Adb00010010010	(	adb00010010010,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m110111_0	),
Adb00010010011	(	adb00010010011,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m110111_0	),
Adb00010010100	(	adb00010010100,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m110111_0	),
Adb00010010101	(	adb00010010101,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m110111_0	),
Adb00010010110	(	adb00010010110,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m110111_0	),
Adb00010010111	(	adb00010010111,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m110111_0	),
Adb00010011000	(	adb00010011000,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m110111_0	),
Adb00010011001	(	adb00010011001,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m110111_0	),
Adb00010011010	(	adb00010011010,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m110111_0	),
Adb00010011011	(	adb00010011011,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m110111_0	),
Adb00010011100	(	adb00010011100,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m110111_0	),
Adb00010011101	(	adb00010011101,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m110111_0	),
Adb00010011110	(	adb00010011110,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m110111_0	),
Adb00010011111	(	adb00010011111,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m110111_0	),
Adb00010100000	(	adb00010100000,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m110111_0	),
Adb00010100001	(	adb00010100001,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m110111_0	),
Adb00010100010	(	adb00010100010,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m110111_0	),
Adb00010100011	(	adb00010100011,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m110111_0	),
Adb00010100100	(	adb00010100100,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m110111_0	),
Adb00010100101	(	adb00010100101,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m110111_0	),
Adb00010100110	(	adb00010100110,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m110111_0	),
Adb00010100111	(	adb00010100111,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m110111_0	),
Adb00010101000	(	adb00010101000,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m110111_0	),
Adb00010101001	(	adb00010101001,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m110111_0	),
Adb00010101010	(	adb00010101010,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m110111_0	),
Adb00010101011	(	adb00010101011,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m110111_0	),
Adb00010101100	(	adb00010101100,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m110111_0	),
Adb00010101101	(	adb00010101101,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m110111_0	),
Adb00010101110	(	adb00010101110,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m110111_0	),
Adb00010101111	(	adb00010101111,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m110111_0	),
Adb00010110000	(	adb00010110000,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m110111_0	),
Adb00010110001	(	adb00010110001,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m110111_0	),
Adb00010110010	(	adb00010110010,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m110111_0	),
Adb00010110011	(	adb00010110011,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m110111_0	),
Adb00010110100	(	adb00010110100,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m110111_0	),
Adb00010110101	(	adb00010110101,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m110111_0	),
Adb00010110110	(	adb00010110110,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m110111_0	),
Adb00010110111	(	adb00010110111,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m110111_0	),
Adb00010111000	(	adb00010111000,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m110111_0	),
Adb00010111001	(	adb00010111001,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m110111_0	),
Adb00010111010	(	adb00010111010,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m110111_0	),
Adb00010111011	(	adb00010111011,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m110111_0	),
Adb00010111100	(	adb00010111100,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m110111_0	),
Adb00010111101	(	adb00010111101,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m110111_0	),
Adb00010111110	(	adb00010111110,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m110111_0	),
Adb00010111111	(	adb00010111111,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m110111_0	),
Adb00011000000	(	adb00011000000,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m110111_0	),
Adb00011000001	(	adb00011000001,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m110111_0	),
Adb00011000010	(	adb00011000010,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m110111_0	),
Adb00011000011	(	adb00011000011,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m110111_0	),
Adb00011000100	(	adb00011000100,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m110111_0	),
Adb00011000101	(	adb00011000101,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m110111_0	),
Adb00011000110	(	adb00011000110,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m110111_0	),
Adb00011000111	(	adb00011000111,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m110111_0	),
Adb00011001000	(	adb00011001000,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m110111_0	),
Adb00011001001	(	adb00011001001,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m110111_0	),
Adb00011001010	(	adb00011001010,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m110111_0	),
Adb00011001011	(	adb00011001011,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m110111_0	),
Adb00011001100	(	adb00011001100,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m110111_0	),
Adb00011001101	(	adb00011001101,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m110111_0	),
Adb00011001110	(	adb00011001110,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m110111_0	),
Adb00011001111	(	adb00011001111,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m110111_0	),
Adb00011010000	(	adb00011010000,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m110111_0	),
Adb00011010001	(	adb00011010001,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m110111_0	),
Adb00011010010	(	adb00011010010,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m110111_0	),
Adb00011010011	(	adb00011010011,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m110111_0	),
Adb00011010100	(	adb00011010100,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m110111_0	),
Adb00011010101	(	adb00011010101,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m110111_0	),
Adb00011010110	(	adb00011010110,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m110111_0	),
Adb00011010111	(	adb00011010111,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m110111_0	),
Adb00011011000	(	adb00011011000,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m110111_0	),
Adb00011011001	(	adb00011011001,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m110111_0	),
Adb00011011010	(	adb00011011010,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m110111_0	),
Adb00011011011	(	adb00011011011,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m110111_0	),
Adb00011011100	(	adb00011011100,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m110111_0	),
Adb00011011101	(	adb00011011101,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m110111_0	),
Adb00011011110	(	adb00011011110,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m110111_0	),
Adb00011011111	(	adb00011011111,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m110111_0	),
Adb00011100000	(	adb00011100000,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m110111_0	),
Adb00011100001	(	adb00011100001,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m110111_0	),
Adb00011100010	(	adb00011100010,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m110111_0	),
Adb00011100011	(	adb00011100011,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m110111_0	),
Adb00011100100	(	adb00011100100,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m110111_0	),
Adb00011100101	(	adb00011100101,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m110111_0	),
Adb00011100110	(	adb00011100110,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m110111_0	),
Adb00011100111	(	adb00011100111,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m110111_0	),
Adb00011101000	(	adb00011101000,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m110111_0	),
Adb00011101001	(	adb00011101001,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m110111_0	),
Adb00011101010	(	adb00011101010,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m110111_0	),
Adb00011101011	(	adb00011101011,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m110111_0	),
Adb00011101100	(	adb00011101100,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m110111_0	),
Adb00011101101	(	adb00011101101,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m110111_0	),
Adb00011101110	(	adb00011101110,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m110111_0	),
Adb00011101111	(	adb00011101111,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m110111_0	),
Adb00011110000	(	adb00011110000,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m110111_0	),
Adb00011110001	(	adb00011110001,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m110111_0	),
Adb00011110010	(	adb00011110010,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m110111_0	),
Adb00011110011	(	adb00011110011,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m110111_0	),
Adb00011110100	(	adb00011110100,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m110111_0	),
Adb00011110101	(	adb00011110101,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m110111_0	),
Adb00011110110	(	adb00011110110,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m110111_0	),
Adb00011110111	(	adb00011110111,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m110111_0	),
Adb00011111000	(	adb00011111000,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m110111_0	),
Adb00011111001	(	adb00011111001,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m110111_0	),
Adb00011111010	(	adb00011111010,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m110111_0	),
Adb00011111011	(	adb00011111011,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m110111_0	),
Adb00011111100	(	adb00011111100,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m110111_0	),
Adb00011111101	(	adb00011111101,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m110111_0	),
Adb00011111110	(	adb00011111110,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m110111_0	),
Adb00011111111	(	adb00011111111,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m110111_0	),
Adb00100000000	(	adb00100000000,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m101111_0	),
Adb00100000001	(	adb00100000001,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m101111_0	),
Adb00100000010	(	adb00100000010,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m101111_0	),
Adb00100000011	(	adb00100000011,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m101111_0	),
Adb00100000100	(	adb00100000100,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m101111_0	),
Adb00100000101	(	adb00100000101,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m101111_0	),
Adb00100000110	(	adb00100000110,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m101111_0	),
Adb00100000111	(	adb00100000111,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m101111_0	),
Adb00100001000	(	adb00100001000,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m101111_0	),
Adb00100001001	(	adb00100001001,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m101111_0	),
Adb00100001010	(	adb00100001010,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m101111_0	),
Adb00100001011	(	adb00100001011,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m101111_0	),
Adb00100001100	(	adb00100001100,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m101111_0	),
Adb00100001101	(	adb00100001101,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m101111_0	),
Adb00100001110	(	adb00100001110,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m101111_0	),
Adb00100001111	(	adb00100001111,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m101111_0	),
Adb00100010000	(	adb00100010000,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m101111_0	),
Adb00100010001	(	adb00100010001,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m101111_0	),
Adb00100010010	(	adb00100010010,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m101111_0	),
Adb00100010011	(	adb00100010011,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m101111_0	),
Adb00100010100	(	adb00100010100,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m101111_0	),
Adb00100010101	(	adb00100010101,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m101111_0	),
Adb00100010110	(	adb00100010110,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m101111_0	),
Adb00100010111	(	adb00100010111,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m101111_0	),
Adb00100011000	(	adb00100011000,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m101111_0	),
Adb00100011001	(	adb00100011001,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m101111_0	),
Adb00100011010	(	adb00100011010,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m101111_0	),
Adb00100011011	(	adb00100011011,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m101111_0	),
Adb00100011100	(	adb00100011100,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m101111_0	),
Adb00100011101	(	adb00100011101,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m101111_0	),
Adb00100011110	(	adb00100011110,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m101111_0	),
Adb00100011111	(	adb00100011111,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m101111_0	),
Adb00100100000	(	adb00100100000,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m101111_0	),
Adb00100100001	(	adb00100100001,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m101111_0	),
Adb00100100010	(	adb00100100010,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m101111_0	),
Adb00100100011	(	adb00100100011,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m101111_0	),
Adb00100100100	(	adb00100100100,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m101111_0	),
Adb00100100101	(	adb00100100101,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m101111_0	),
Adb00100100110	(	adb00100100110,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m101111_0	),
Adb00100100111	(	adb00100100111,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m101111_0	),
Adb00100101000	(	adb00100101000,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m101111_0	),
Adb00100101001	(	adb00100101001,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m101111_0	),
Adb00100101010	(	adb00100101010,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m101111_0	),
Adb00100101011	(	adb00100101011,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m101111_0	),
Adb00100101100	(	adb00100101100,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m101111_0	),
Adb00100101101	(	adb00100101101,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m101111_0	),
Adb00100101110	(	adb00100101110,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m101111_0	),
Adb00100101111	(	adb00100101111,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m101111_0	),
Adb00100110000	(	adb00100110000,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m101111_0	),
Adb00100110001	(	adb00100110001,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m101111_0	),
Adb00100110010	(	adb00100110010,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m101111_0	),
Adb00100110011	(	adb00100110011,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m101111_0	),
Adb00100110100	(	adb00100110100,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m101111_0	),
Adb00100110101	(	adb00100110101,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m101111_0	),
Adb00100110110	(	adb00100110110,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m101111_0	),
Adb00100110111	(	adb00100110111,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m101111_0	),
Adb00100111000	(	adb00100111000,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m101111_0	),
Adb00100111001	(	adb00100111001,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m101111_0	),
Adb00100111010	(	adb00100111010,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m101111_0	),
Adb00100111011	(	adb00100111011,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m101111_0	),
Adb00100111100	(	adb00100111100,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m101111_0	),
Adb00100111101	(	adb00100111101,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m101111_0	),
Adb00100111110	(	adb00100111110,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m101111_0	),
Adb00100111111	(	adb00100111111,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m101111_0	),
Adb00101000000	(	adb00101000000,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m101111_0	),
Adb00101000001	(	adb00101000001,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m101111_0	),
Adb00101000010	(	adb00101000010,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m101111_0	),
Adb00101000011	(	adb00101000011,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m101111_0	),
Adb00101000100	(	adb00101000100,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m101111_0	),
Adb00101000101	(	adb00101000101,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m101111_0	),
Adb00101000110	(	adb00101000110,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m101111_0	),
Adb00101000111	(	adb00101000111,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m101111_0	),
Adb00101001000	(	adb00101001000,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m101111_0	),
Adb00101001001	(	adb00101001001,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m101111_0	),
Adb00101001010	(	adb00101001010,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m101111_0	),
Adb00101001011	(	adb00101001011,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m101111_0	),
Adb00101001100	(	adb00101001100,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m101111_0	),
Adb00101001101	(	adb00101001101,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m101111_0	),
Adb00101001110	(	adb00101001110,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m101111_0	),
Adb00101001111	(	adb00101001111,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m101111_0	),
Adb00101010000	(	adb00101010000,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m101111_0	),
Adb00101010001	(	adb00101010001,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m101111_0	),
Adb00101010010	(	adb00101010010,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m101111_0	),
Adb00101010011	(	adb00101010011,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m101111_0	),
Adb00101010100	(	adb00101010100,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m101111_0	),
Adb00101010101	(	adb00101010101,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m101111_0	),
Adb00101010110	(	adb00101010110,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m101111_0	),
Adb00101010111	(	adb00101010111,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m101111_0	),
Adb00101011000	(	adb00101011000,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m101111_0	),
Adb00101011001	(	adb00101011001,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m101111_0	),
Adb00101011010	(	adb00101011010,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m101111_0	),
Adb00101011011	(	adb00101011011,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m101111_0	),
Adb00101011100	(	adb00101011100,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m101111_0	),
Adb00101011101	(	adb00101011101,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m101111_0	),
Adb00101011110	(	adb00101011110,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m101111_0	),
Adb00101011111	(	adb00101011111,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m101111_0	),
Adb00101100000	(	adb00101100000,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m101111_0	),
Adb00101100001	(	adb00101100001,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m101111_0	),
Adb00101100010	(	adb00101100010,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m101111_0	),
Adb00101100011	(	adb00101100011,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m101111_0	),
Adb00101100100	(	adb00101100100,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m101111_0	),
Adb00101100101	(	adb00101100101,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m101111_0	),
Adb00101100110	(	adb00101100110,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m101111_0	),
Adb00101100111	(	adb00101100111,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m101111_0	),
Adb00101101000	(	adb00101101000,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m101111_0	),
Adb00101101001	(	adb00101101001,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m101111_0	),
Adb00101101010	(	adb00101101010,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m101111_0	),
Adb00101101011	(	adb00101101011,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m101111_0	),
Adb00101101100	(	adb00101101100,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m101111_0	),
Adb00101101101	(	adb00101101101,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m101111_0	),
Adb00101101110	(	adb00101101110,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m101111_0	),
Adb00101101111	(	adb00101101111,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m101111_0	),
Adb00101110000	(	adb00101110000,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m101111_0	),
Adb00101110001	(	adb00101110001,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m101111_0	),
Adb00101110010	(	adb00101110010,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m101111_0	),
Adb00101110011	(	adb00101110011,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m101111_0	),
Adb00101110100	(	adb00101110100,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m101111_0	),
Adb00101110101	(	adb00101110101,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m101111_0	),
Adb00101110110	(	adb00101110110,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m101111_0	),
Adb00101110111	(	adb00101110111,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m101111_0	),
Adb00101111000	(	adb00101111000,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m101111_0	),
Adb00101111001	(	adb00101111001,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m101111_0	),
Adb00101111010	(	adb00101111010,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m101111_0	),
Adb00101111011	(	adb00101111011,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m101111_0	),
Adb00101111100	(	adb00101111100,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m101111_0	),
Adb00101111101	(	adb00101111101,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m101111_0	),
Adb00101111110	(	adb00101111110,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m101111_0	),
Adb00101111111	(	adb00101111111,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m101111_0	),
Adb00110000000	(	adb00110000000,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m100111_0	),
Adb00110000001	(	adb00110000001,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m100111_0	),
Adb00110000010	(	adb00110000010,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m100111_0	),
Adb00110000011	(	adb00110000011,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m100111_0	),
Adb00110000100	(	adb00110000100,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m100111_0	),
Adb00110000101	(	adb00110000101,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m100111_0	),
Adb00110000110	(	adb00110000110,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m100111_0	),
Adb00110000111	(	adb00110000111,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m100111_0	),
Adb00110001000	(	adb00110001000,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m100111_0	),
Adb00110001001	(	adb00110001001,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m100111_0	),
Adb00110001010	(	adb00110001010,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m100111_0	),
Adb00110001011	(	adb00110001011,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m100111_0	),
Adb00110001100	(	adb00110001100,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m100111_0	),
Adb00110001101	(	adb00110001101,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m100111_0	),
Adb00110001110	(	adb00110001110,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m100111_0	),
Adb00110001111	(	adb00110001111,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m100111_0	),
Adb00110010000	(	adb00110010000,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m100111_0	),
Adb00110010001	(	adb00110010001,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m100111_0	),
Adb00110010010	(	adb00110010010,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m100111_0	),
Adb00110010011	(	adb00110010011,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m100111_0	),
Adb00110010100	(	adb00110010100,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m100111_0	),
Adb00110010101	(	adb00110010101,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m100111_0	),
Adb00110010110	(	adb00110010110,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m100111_0	),
Adb00110010111	(	adb00110010111,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m100111_0	),
Adb00110011000	(	adb00110011000,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m100111_0	),
Adb00110011001	(	adb00110011001,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m100111_0	),
Adb00110011010	(	adb00110011010,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m100111_0	),
Adb00110011011	(	adb00110011011,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m100111_0	),
Adb00110011100	(	adb00110011100,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m100111_0	),
Adb00110011101	(	adb00110011101,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m100111_0	),
Adb00110011110	(	adb00110011110,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m100111_0	),
Adb00110011111	(	adb00110011111,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m100111_0	),
Adb00110100000	(	adb00110100000,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m100111_0	),
Adb00110100001	(	adb00110100001,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m100111_0	),
Adb00110100010	(	adb00110100010,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m100111_0	),
Adb00110100011	(	adb00110100011,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m100111_0	),
Adb00110100100	(	adb00110100100,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m100111_0	),
Adb00110100101	(	adb00110100101,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m100111_0	),
Adb00110100110	(	adb00110100110,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m100111_0	),
Adb00110100111	(	adb00110100111,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m100111_0	),
Adb00110101000	(	adb00110101000,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m100111_0	),
Adb00110101001	(	adb00110101001,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m100111_0	),
Adb00110101010	(	adb00110101010,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m100111_0	),
Adb00110101011	(	adb00110101011,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m100111_0	),
Adb00110101100	(	adb00110101100,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m100111_0	),
Adb00110101101	(	adb00110101101,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m100111_0	),
Adb00110101110	(	adb00110101110,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m100111_0	),
Adb00110101111	(	adb00110101111,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m100111_0	),
Adb00110110000	(	adb00110110000,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m100111_0	),
Adb00110110001	(	adb00110110001,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m100111_0	),
Adb00110110010	(	adb00110110010,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m100111_0	),
Adb00110110011	(	adb00110110011,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m100111_0	),
Adb00110110100	(	adb00110110100,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m100111_0	),
Adb00110110101	(	adb00110110101,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m100111_0	),
Adb00110110110	(	adb00110110110,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m100111_0	),
Adb00110110111	(	adb00110110111,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m100111_0	),
Adb00110111000	(	adb00110111000,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m100111_0	),
Adb00110111001	(	adb00110111001,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m100111_0	),
Adb00110111010	(	adb00110111010,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m100111_0	),
Adb00110111011	(	adb00110111011,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m100111_0	),
Adb00110111100	(	adb00110111100,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m100111_0	),
Adb00110111101	(	adb00110111101,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m100111_0	),
Adb00110111110	(	adb00110111110,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m100111_0	),
Adb00110111111	(	adb00110111111,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m100111_0	),
Adb00111000000	(	adb00111000000,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m100111_0	),
Adb00111000001	(	adb00111000001,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m100111_0	),
Adb00111000010	(	adb00111000010,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m100111_0	),
Adb00111000011	(	adb00111000011,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m100111_0	),
Adb00111000100	(	adb00111000100,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m100111_0	),
Adb00111000101	(	adb00111000101,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m100111_0	),
Adb00111000110	(	adb00111000110,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m100111_0	),
Adb00111000111	(	adb00111000111,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m100111_0	),
Adb00111001000	(	adb00111001000,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m100111_0	),
Adb00111001001	(	adb00111001001,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m100111_0	),
Adb00111001010	(	adb00111001010,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m100111_0	),
Adb00111001011	(	adb00111001011,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m100111_0	),
Adb00111001100	(	adb00111001100,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m100111_0	),
Adb00111001101	(	adb00111001101,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m100111_0	),
Adb00111001110	(	adb00111001110,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m100111_0	),
Adb00111001111	(	adb00111001111,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m100111_0	),
Adb00111010000	(	adb00111010000,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m100111_0	),
Adb00111010001	(	adb00111010001,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m100111_0	),
Adb00111010010	(	adb00111010010,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m100111_0	),
Adb00111010011	(	adb00111010011,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m100111_0	),
Adb00111010100	(	adb00111010100,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m100111_0	),
Adb00111010101	(	adb00111010101,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m100111_0	),
Adb00111010110	(	adb00111010110,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m100111_0	),
Adb00111010111	(	adb00111010111,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m100111_0	),
Adb00111011000	(	adb00111011000,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m100111_0	),
Adb00111011001	(	adb00111011001,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m100111_0	),
Adb00111011010	(	adb00111011010,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m100111_0	),
Adb00111011011	(	adb00111011011,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m100111_0	),
Adb00111011100	(	adb00111011100,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m100111_0	),
Adb00111011101	(	adb00111011101,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m100111_0	),
Adb00111011110	(	adb00111011110,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m100111_0	),
Adb00111011111	(	adb00111011111,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m100111_0	),
Adb00111100000	(	adb00111100000,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m100111_0	),
Adb00111100001	(	adb00111100001,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m100111_0	),
Adb00111100010	(	adb00111100010,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m100111_0	),
Adb00111100011	(	adb00111100011,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m100111_0	),
Adb00111100100	(	adb00111100100,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m100111_0	),
Adb00111100101	(	adb00111100101,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m100111_0	),
Adb00111100110	(	adb00111100110,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m100111_0	),
Adb00111100111	(	adb00111100111,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m100111_0	),
Adb00111101000	(	adb00111101000,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m100111_0	),
Adb00111101001	(	adb00111101001,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m100111_0	),
Adb00111101010	(	adb00111101010,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m100111_0	),
Adb00111101011	(	adb00111101011,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m100111_0	),
Adb00111101100	(	adb00111101100,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m100111_0	),
Adb00111101101	(	adb00111101101,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m100111_0	),
Adb00111101110	(	adb00111101110,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m100111_0	),
Adb00111101111	(	adb00111101111,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m100111_0	),
Adb00111110000	(	adb00111110000,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m100111_0	),
Adb00111110001	(	adb00111110001,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m100111_0	),
Adb00111110010	(	adb00111110010,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m100111_0	),
Adb00111110011	(	adb00111110011,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m100111_0	),
Adb00111110100	(	adb00111110100,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m100111_0	),
Adb00111110101	(	adb00111110101,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m100111_0	),
Adb00111110110	(	adb00111110110,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m100111_0	),
Adb00111110111	(	adb00111110111,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m100111_0	),
Adb00111111000	(	adb00111111000,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m100111_0	),
Adb00111111001	(	adb00111111001,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m100111_0	),
Adb00111111010	(	adb00111111010,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m100111_0	),
Adb00111111011	(	adb00111111011,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m100111_0	),
Adb00111111100	(	adb00111111100,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m100111_0	),
Adb00111111101	(	adb00111111101,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m100111_0	),
Adb00111111110	(	adb00111111110,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m100111_0	),
Adb00111111111	(	adb00111111111,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m100111_0	),
Adb01000000000	(	adb01000000000,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m011111_0	),
Adb01000000001	(	adb01000000001,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m011111_0	),
Adb01000000010	(	adb01000000010,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m011111_0	),
Adb01000000011	(	adb01000000011,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m011111_0	),
Adb01000000100	(	adb01000000100,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m011111_0	),
Adb01000000101	(	adb01000000101,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m011111_0	),
Adb01000000110	(	adb01000000110,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m011111_0	),
Adb01000000111	(	adb01000000111,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m011111_0	),
Adb01000001000	(	adb01000001000,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m011111_0	),
Adb01000001001	(	adb01000001001,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m011111_0	),
Adb01000001010	(	adb01000001010,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m011111_0	),
Adb01000001011	(	adb01000001011,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m011111_0	),
Adb01000001100	(	adb01000001100,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m011111_0	),
Adb01000001101	(	adb01000001101,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m011111_0	),
Adb01000001110	(	adb01000001110,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m011111_0	),
Adb01000001111	(	adb01000001111,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m011111_0	),
Adb01000010000	(	adb01000010000,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m011111_0	),
Adb01000010001	(	adb01000010001,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m011111_0	),
Adb01000010010	(	adb01000010010,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m011111_0	),
Adb01000010011	(	adb01000010011,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m011111_0	),
Adb01000010100	(	adb01000010100,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m011111_0	),
Adb01000010101	(	adb01000010101,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m011111_0	),
Adb01000010110	(	adb01000010110,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m011111_0	),
Adb01000010111	(	adb01000010111,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m011111_0	),
Adb01000011000	(	adb01000011000,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m011111_0	),
Adb01000011001	(	adb01000011001,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m011111_0	),
Adb01000011010	(	adb01000011010,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m011111_0	),
Adb01000011011	(	adb01000011011,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m011111_0	),
Adb01000011100	(	adb01000011100,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m011111_0	),
Adb01000011101	(	adb01000011101,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m011111_0	),
Adb01000011110	(	adb01000011110,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m011111_0	),
Adb01000011111	(	adb01000011111,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m011111_0	),
Adb01000100000	(	adb01000100000,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m011111_0	),
Adb01000100001	(	adb01000100001,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m011111_0	),
Adb01000100010	(	adb01000100010,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m011111_0	),
Adb01000100011	(	adb01000100011,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m011111_0	),
Adb01000100100	(	adb01000100100,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m011111_0	),
Adb01000100101	(	adb01000100101,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m011111_0	),
Adb01000100110	(	adb01000100110,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m011111_0	),
Adb01000100111	(	adb01000100111,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m011111_0	),
Adb01000101000	(	adb01000101000,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m011111_0	),
Adb01000101001	(	adb01000101001,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m011111_0	),
Adb01000101010	(	adb01000101010,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m011111_0	),
Adb01000101011	(	adb01000101011,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m011111_0	),
Adb01000101100	(	adb01000101100,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m011111_0	),
Adb01000101101	(	adb01000101101,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m011111_0	),
Adb01000101110	(	adb01000101110,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m011111_0	),
Adb01000101111	(	adb01000101111,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m011111_0	),
Adb01000110000	(	adb01000110000,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m011111_0	),
Adb01000110001	(	adb01000110001,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m011111_0	),
Adb01000110010	(	adb01000110010,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m011111_0	),
Adb01000110011	(	adb01000110011,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m011111_0	),
Adb01000110100	(	adb01000110100,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m011111_0	),
Adb01000110101	(	adb01000110101,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m011111_0	),
Adb01000110110	(	adb01000110110,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m011111_0	),
Adb01000110111	(	adb01000110111,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m011111_0	),
Adb01000111000	(	adb01000111000,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m011111_0	),
Adb01000111001	(	adb01000111001,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m011111_0	),
Adb01000111010	(	adb01000111010,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m011111_0	),
Adb01000111011	(	adb01000111011,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m011111_0	),
Adb01000111100	(	adb01000111100,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m011111_0	),
Adb01000111101	(	adb01000111101,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m011111_0	),
Adb01000111110	(	adb01000111110,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m011111_0	),
Adb01000111111	(	adb01000111111,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m011111_0	),
Adb01001000000	(	adb01001000000,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m011111_0	),
Adb01001000001	(	adb01001000001,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m011111_0	),
Adb01001000010	(	adb01001000010,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m011111_0	),
Adb01001000011	(	adb01001000011,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m011111_0	),
Adb01001000100	(	adb01001000100,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m011111_0	),
Adb01001000101	(	adb01001000101,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m011111_0	),
Adb01001000110	(	adb01001000110,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m011111_0	),
Adb01001000111	(	adb01001000111,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m011111_0	),
Adb01001001000	(	adb01001001000,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m011111_0	),
Adb01001001001	(	adb01001001001,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m011111_0	),
Adb01001001010	(	adb01001001010,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m011111_0	),
Adb01001001011	(	adb01001001011,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m011111_0	),
Adb01001001100	(	adb01001001100,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m011111_0	),
Adb01001001101	(	adb01001001101,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m011111_0	),
Adb01001001110	(	adb01001001110,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m011111_0	),
Adb01001001111	(	adb01001001111,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m011111_0	),
Adb01001010000	(	adb01001010000,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m011111_0	),
Adb01001010001	(	adb01001010001,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m011111_0	),
Adb01001010010	(	adb01001010010,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m011111_0	),
Adb01001010011	(	adb01001010011,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m011111_0	),
Adb01001010100	(	adb01001010100,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m011111_0	),
Adb01001010101	(	adb01001010101,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m011111_0	),
Adb01001010110	(	adb01001010110,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m011111_0	),
Adb01001010111	(	adb01001010111,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m011111_0	),
Adb01001011000	(	adb01001011000,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m011111_0	),
Adb01001011001	(	adb01001011001,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m011111_0	),
Adb01001011010	(	adb01001011010,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m011111_0	),
Adb01001011011	(	adb01001011011,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m011111_0	),
Adb01001011100	(	adb01001011100,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m011111_0	),
Adb01001011101	(	adb01001011101,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m011111_0	),
Adb01001011110	(	adb01001011110,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m011111_0	),
Adb01001011111	(	adb01001011111,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m011111_0	),
Adb01001100000	(	adb01001100000,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m011111_0	),
Adb01001100001	(	adb01001100001,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m011111_0	),
Adb01001100010	(	adb01001100010,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m011111_0	),
Adb01001100011	(	adb01001100011,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m011111_0	),
Adb01001100100	(	adb01001100100,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m011111_0	),
Adb01001100101	(	adb01001100101,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m011111_0	),
Adb01001100110	(	adb01001100110,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m011111_0	),
Adb01001100111	(	adb01001100111,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m011111_0	),
Adb01001101000	(	adb01001101000,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m011111_0	),
Adb01001101001	(	adb01001101001,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m011111_0	),
Adb01001101010	(	adb01001101010,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m011111_0	),
Adb01001101011	(	adb01001101011,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m011111_0	),
Adb01001101100	(	adb01001101100,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m011111_0	),
Adb01001101101	(	adb01001101101,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m011111_0	),
Adb01001101110	(	adb01001101110,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m011111_0	),
Adb01001101111	(	adb01001101111,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m011111_0	),
Adb01001110000	(	adb01001110000,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m011111_0	),
Adb01001110001	(	adb01001110001,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m011111_0	),
Adb01001110010	(	adb01001110010,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m011111_0	),
Adb01001110011	(	adb01001110011,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m011111_0	),
Adb01001110100	(	adb01001110100,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m011111_0	),
Adb01001110101	(	adb01001110101,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m011111_0	),
Adb01001110110	(	adb01001110110,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m011111_0	),
Adb01001110111	(	adb01001110111,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m011111_0	),
Adb01001111000	(	adb01001111000,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m011111_0	),
Adb01001111001	(	adb01001111001,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m011111_0	),
Adb01001111010	(	adb01001111010,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m011111_0	),
Adb01001111011	(	adb01001111011,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m011111_0	),
Adb01001111100	(	adb01001111100,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m011111_0	),
Adb01001111101	(	adb01001111101,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m011111_0	),
Adb01001111110	(	adb01001111110,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m011111_0	),
Adb01001111111	(	adb01001111111,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m011111_0	),
Adb01010000000	(	adb01010000000,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m010111_0	),
Adb01010000001	(	adb01010000001,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m010111_0	),
Adb01010000010	(	adb01010000010,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m010111_0	),
Adb01010000011	(	adb01010000011,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m010111_0	),
Adb01010000100	(	adb01010000100,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m010111_0	),
Adb01010000101	(	adb01010000101,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m010111_0	),
Adb01010000110	(	adb01010000110,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m010111_0	),
Adb01010000111	(	adb01010000111,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m010111_0	),
Adb01010001000	(	adb01010001000,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m010111_0	),
Adb01010001001	(	adb01010001001,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m010111_0	),
Adb01010001010	(	adb01010001010,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m010111_0	),
Adb01010001011	(	adb01010001011,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m010111_0	),
Adb01010001100	(	adb01010001100,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m010111_0	),
Adb01010001101	(	adb01010001101,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m010111_0	),
Adb01010001110	(	adb01010001110,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m010111_0	),
Adb01010001111	(	adb01010001111,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m010111_0	),
Adb01010010000	(	adb01010010000,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m010111_0	),
Adb01010010001	(	adb01010010001,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m010111_0	),
Adb01010010010	(	adb01010010010,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m010111_0	),
Adb01010010011	(	adb01010010011,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m010111_0	),
Adb01010010100	(	adb01010010100,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m010111_0	),
Adb01010010101	(	adb01010010101,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m010111_0	),
Adb01010010110	(	adb01010010110,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m010111_0	),
Adb01010010111	(	adb01010010111,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m010111_0	),
Adb01010011000	(	adb01010011000,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m010111_0	),
Adb01010011001	(	adb01010011001,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m010111_0	),
Adb01010011010	(	adb01010011010,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m010111_0	),
Adb01010011011	(	adb01010011011,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m010111_0	),
Adb01010011100	(	adb01010011100,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m010111_0	),
Adb01010011101	(	adb01010011101,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m010111_0	),
Adb01010011110	(	adb01010011110,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m010111_0	),
Adb01010011111	(	adb01010011111,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m010111_0	),
Adb01010100000	(	adb01010100000,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m010111_0	),
Adb01010100001	(	adb01010100001,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m010111_0	),
Adb01010100010	(	adb01010100010,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m010111_0	),
Adb01010100011	(	adb01010100011,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m010111_0	),
Adb01010100100	(	adb01010100100,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m010111_0	),
Adb01010100101	(	adb01010100101,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m010111_0	),
Adb01010100110	(	adb01010100110,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m010111_0	),
Adb01010100111	(	adb01010100111,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m010111_0	),
Adb01010101000	(	adb01010101000,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m010111_0	),
Adb01010101001	(	adb01010101001,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m010111_0	),
Adb01010101010	(	adb01010101010,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m010111_0	),
Adb01010101011	(	adb01010101011,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m010111_0	),
Adb01010101100	(	adb01010101100,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m010111_0	),
Adb01010101101	(	adb01010101101,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m010111_0	),
Adb01010101110	(	adb01010101110,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m010111_0	),
Adb01010101111	(	adb01010101111,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m010111_0	),
Adb01010110000	(	adb01010110000,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m010111_0	),
Adb01010110001	(	adb01010110001,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m010111_0	),
Adb01010110010	(	adb01010110010,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m010111_0	),
Adb01010110011	(	adb01010110011,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m010111_0	),
Adb01010110100	(	adb01010110100,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m010111_0	),
Adb01010110101	(	adb01010110101,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m010111_0	),
Adb01010110110	(	adb01010110110,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m010111_0	),
Adb01010110111	(	adb01010110111,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m010111_0	),
Adb01010111000	(	adb01010111000,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m010111_0	),
Adb01010111001	(	adb01010111001,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m010111_0	),
Adb01010111010	(	adb01010111010,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m010111_0	),
Adb01010111011	(	adb01010111011,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m010111_0	),
Adb01010111100	(	adb01010111100,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m010111_0	),
Adb01010111101	(	adb01010111101,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m010111_0	),
Adb01010111110	(	adb01010111110,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m010111_0	),
Adb01010111111	(	adb01010111111,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m010111_0	),
Adb01011000000	(	adb01011000000,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m010111_0	),
Adb01011000001	(	adb01011000001,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m010111_0	),
Adb01011000010	(	adb01011000010,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m010111_0	),
Adb01011000011	(	adb01011000011,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m010111_0	),
Adb01011000100	(	adb01011000100,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m010111_0	),
Adb01011000101	(	adb01011000101,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m010111_0	),
Adb01011000110	(	adb01011000110,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m010111_0	),
Adb01011000111	(	adb01011000111,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m010111_0	),
Adb01011001000	(	adb01011001000,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m010111_0	),
Adb01011001001	(	adb01011001001,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m010111_0	),
Adb01011001010	(	adb01011001010,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m010111_0	),
Adb01011001011	(	adb01011001011,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m010111_0	),
Adb01011001100	(	adb01011001100,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m010111_0	),
Adb01011001101	(	adb01011001101,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m010111_0	),
Adb01011001110	(	adb01011001110,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m010111_0	),
Adb01011001111	(	adb01011001111,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m010111_0	),
Adb01011010000	(	adb01011010000,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m010111_0	),
Adb01011010001	(	adb01011010001,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m010111_0	),
Adb01011010010	(	adb01011010010,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m010111_0	),
Adb01011010011	(	adb01011010011,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m010111_0	),
Adb01011010100	(	adb01011010100,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m010111_0	),
Adb01011010101	(	adb01011010101,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m010111_0	),
Adb01011010110	(	adb01011010110,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m010111_0	),
Adb01011010111	(	adb01011010111,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m010111_0	),
Adb01011011000	(	adb01011011000,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m010111_0	),
Adb01011011001	(	adb01011011001,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m010111_0	),
Adb01011011010	(	adb01011011010,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m010111_0	),
Adb01011011011	(	adb01011011011,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m010111_0	),
Adb01011011100	(	adb01011011100,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m010111_0	),
Adb01011011101	(	adb01011011101,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m010111_0	),
Adb01011011110	(	adb01011011110,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m010111_0	),
Adb01011011111	(	adb01011011111,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m010111_0	),
Adb01011100000	(	adb01011100000,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m010111_0	),
Adb01011100001	(	adb01011100001,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m010111_0	),
Adb01011100010	(	adb01011100010,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m010111_0	),
Adb01011100011	(	adb01011100011,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m010111_0	),
Adb01011100100	(	adb01011100100,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m010111_0	),
Adb01011100101	(	adb01011100101,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m010111_0	),
Adb01011100110	(	adb01011100110,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m010111_0	),
Adb01011100111	(	adb01011100111,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m010111_0	),
Adb01011101000	(	adb01011101000,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m010111_0	),
Adb01011101001	(	adb01011101001,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m010111_0	),
Adb01011101010	(	adb01011101010,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m010111_0	),
Adb01011101011	(	adb01011101011,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m010111_0	),
Adb01011101100	(	adb01011101100,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m010111_0	),
Adb01011101101	(	adb01011101101,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m010111_0	),
Adb01011101110	(	adb01011101110,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m010111_0	),
Adb01011101111	(	adb01011101111,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m010111_0	),
Adb01011110000	(	adb01011110000,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m010111_0	),
Adb01011110001	(	adb01011110001,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m010111_0	),
Adb01011110010	(	adb01011110010,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m010111_0	),
Adb01011110011	(	adb01011110011,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m010111_0	),
Adb01011110100	(	adb01011110100,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m010111_0	),
Adb01011110101	(	adb01011110101,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m010111_0	),
Adb01011110110	(	adb01011110110,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m010111_0	),
Adb01011110111	(	adb01011110111,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m010111_0	),
Adb01011111000	(	adb01011111000,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m010111_0	),
Adb01011111001	(	adb01011111001,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m010111_0	),
Adb01011111010	(	adb01011111010,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m010111_0	),
Adb01011111011	(	adb01011111011,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m010111_0	),
Adb01011111100	(	adb01011111100,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m010111_0	),
Adb01011111101	(	adb01011111101,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m010111_0	),
Adb01011111110	(	adb01011111110,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m010111_0	),
Adb01011111111	(	adb01011111111,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m010111_0	),
Adb01100000000	(	adb01100000000,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m001111_0	),
Adb01100000001	(	adb01100000001,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m001111_0	),
Adb01100000010	(	adb01100000010,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m001111_0	),
Adb01100000011	(	adb01100000011,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m001111_0	),
Adb01100000100	(	adb01100000100,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m001111_0	),
Adb01100000101	(	adb01100000101,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m001111_0	),
Adb01100000110	(	adb01100000110,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m001111_0	),
Adb01100000111	(	adb01100000111,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m001111_0	),
Adb01100001000	(	adb01100001000,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m001111_0	),
Adb01100001001	(	adb01100001001,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m001111_0	),
Adb01100001010	(	adb01100001010,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m001111_0	),
Adb01100001011	(	adb01100001011,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m001111_0	),
Adb01100001100	(	adb01100001100,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m001111_0	),
Adb01100001101	(	adb01100001101,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m001111_0	),
Adb01100001110	(	adb01100001110,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m001111_0	),
Adb01100001111	(	adb01100001111,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m001111_0	),
Adb01100010000	(	adb01100010000,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m001111_0	),
Adb01100010001	(	adb01100010001,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m001111_0	),
Adb01100010010	(	adb01100010010,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m001111_0	),
Adb01100010011	(	adb01100010011,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m001111_0	),
Adb01100010100	(	adb01100010100,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m001111_0	),
Adb01100010101	(	adb01100010101,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m001111_0	),
Adb01100010110	(	adb01100010110,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m001111_0	),
Adb01100010111	(	adb01100010111,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m001111_0	),
Adb01100011000	(	adb01100011000,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m001111_0	),
Adb01100011001	(	adb01100011001,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m001111_0	),
Adb01100011010	(	adb01100011010,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m001111_0	),
Adb01100011011	(	adb01100011011,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m001111_0	),
Adb01100011100	(	adb01100011100,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m001111_0	),
Adb01100011101	(	adb01100011101,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m001111_0	),
Adb01100011110	(	adb01100011110,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m001111_0	),
Adb01100011111	(	adb01100011111,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m001111_0	),
Adb01100100000	(	adb01100100000,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m001111_0	),
Adb01100100001	(	adb01100100001,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m001111_0	),
Adb01100100010	(	adb01100100010,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m001111_0	),
Adb01100100011	(	adb01100100011,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m001111_0	),
Adb01100100100	(	adb01100100100,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m001111_0	),
Adb01100100101	(	adb01100100101,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m001111_0	),
Adb01100100110	(	adb01100100110,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m001111_0	),
Adb01100100111	(	adb01100100111,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m001111_0	),
Adb01100101000	(	adb01100101000,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m001111_0	),
Adb01100101001	(	adb01100101001,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m001111_0	),
Adb01100101010	(	adb01100101010,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m001111_0	),
Adb01100101011	(	adb01100101011,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m001111_0	),
Adb01100101100	(	adb01100101100,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m001111_0	),
Adb01100101101	(	adb01100101101,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m001111_0	),
Adb01100101110	(	adb01100101110,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m001111_0	),
Adb01100101111	(	adb01100101111,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m001111_0	),
Adb01100110000	(	adb01100110000,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m001111_0	),
Adb01100110001	(	adb01100110001,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m001111_0	),
Adb01100110010	(	adb01100110010,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m001111_0	),
Adb01100110011	(	adb01100110011,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m001111_0	),
Adb01100110100	(	adb01100110100,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m001111_0	),
Adb01100110101	(	adb01100110101,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m001111_0	),
Adb01100110110	(	adb01100110110,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m001111_0	),
Adb01100110111	(	adb01100110111,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m001111_0	),
Adb01100111000	(	adb01100111000,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m001111_0	),
Adb01100111001	(	adb01100111001,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m001111_0	),
Adb01100111010	(	adb01100111010,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m001111_0	),
Adb01100111011	(	adb01100111011,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m001111_0	),
Adb01100111100	(	adb01100111100,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m001111_0	),
Adb01100111101	(	adb01100111101,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m001111_0	),
Adb01100111110	(	adb01100111110,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m001111_0	),
Adb01100111111	(	adb01100111111,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m001111_0	),
Adb01101000000	(	adb01101000000,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m001111_0	),
Adb01101000001	(	adb01101000001,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m001111_0	),
Adb01101000010	(	adb01101000010,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m001111_0	),
Adb01101000011	(	adb01101000011,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m001111_0	),
Adb01101000100	(	adb01101000100,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m001111_0	),
Adb01101000101	(	adb01101000101,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m001111_0	),
Adb01101000110	(	adb01101000110,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m001111_0	),
Adb01101000111	(	adb01101000111,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m001111_0	),
Adb01101001000	(	adb01101001000,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m001111_0	),
Adb01101001001	(	adb01101001001,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m001111_0	),
Adb01101001010	(	adb01101001010,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m001111_0	),
Adb01101001011	(	adb01101001011,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m001111_0	),
Adb01101001100	(	adb01101001100,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m001111_0	),
Adb01101001101	(	adb01101001101,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m001111_0	),
Adb01101001110	(	adb01101001110,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m001111_0	),
Adb01101001111	(	adb01101001111,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m001111_0	),
Adb01101010000	(	adb01101010000,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m001111_0	),
Adb01101010001	(	adb01101010001,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m001111_0	),
Adb01101010010	(	adb01101010010,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m001111_0	),
Adb01101010011	(	adb01101010011,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m001111_0	),
Adb01101010100	(	adb01101010100,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m001111_0	),
Adb01101010101	(	adb01101010101,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m001111_0	),
Adb01101010110	(	adb01101010110,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m001111_0	),
Adb01101010111	(	adb01101010111,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m001111_0	),
Adb01101011000	(	adb01101011000,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m001111_0	),
Adb01101011001	(	adb01101011001,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m001111_0	),
Adb01101011010	(	adb01101011010,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m001111_0	),
Adb01101011011	(	adb01101011011,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m001111_0	),
Adb01101011100	(	adb01101011100,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m001111_0	),
Adb01101011101	(	adb01101011101,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m001111_0	),
Adb01101011110	(	adb01101011110,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m001111_0	),
Adb01101011111	(	adb01101011111,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m001111_0	),
Adb01101100000	(	adb01101100000,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m001111_0	),
Adb01101100001	(	adb01101100001,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m001111_0	),
Adb01101100010	(	adb01101100010,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m001111_0	),
Adb01101100011	(	adb01101100011,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m001111_0	),
Adb01101100100	(	adb01101100100,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m001111_0	),
Adb01101100101	(	adb01101100101,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m001111_0	),
Adb01101100110	(	adb01101100110,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m001111_0	),
Adb01101100111	(	adb01101100111,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m001111_0	),
Adb01101101000	(	adb01101101000,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m001111_0	),
Adb01101101001	(	adb01101101001,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m001111_0	),
Adb01101101010	(	adb01101101010,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m001111_0	),
Adb01101101011	(	adb01101101011,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m001111_0	),
Adb01101101100	(	adb01101101100,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m001111_0	),
Adb01101101101	(	adb01101101101,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m001111_0	),
Adb01101101110	(	adb01101101110,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m001111_0	),
Adb01101101111	(	adb01101101111,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m001111_0	),
Adb01101110000	(	adb01101110000,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m001111_0	),
Adb01101110001	(	adb01101110001,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m001111_0	),
Adb01101110010	(	adb01101110010,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m001111_0	),
Adb01101110011	(	adb01101110011,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m001111_0	),
Adb01101110100	(	adb01101110100,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m001111_0	),
Adb01101110101	(	adb01101110101,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m001111_0	),
Adb01101110110	(	adb01101110110,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m001111_0	),
Adb01101110111	(	adb01101110111,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m001111_0	),
Adb01101111000	(	adb01101111000,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m001111_0	),
Adb01101111001	(	adb01101111001,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m001111_0	),
Adb01101111010	(	adb01101111010,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m001111_0	),
Adb01101111011	(	adb01101111011,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m001111_0	),
Adb01101111100	(	adb01101111100,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m001111_0	),
Adb01101111101	(	adb01101111101,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m001111_0	),
Adb01101111110	(	adb01101111110,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m001111_0	),
Adb01101111111	(	adb01101111111,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m001111_0	),
Adb01110000000	(	adb01110000000,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m000111_0	),
Adb01110000001	(	adb01110000001,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m000111_0	),
Adb01110000010	(	adb01110000010,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m000111_0	),
Adb01110000011	(	adb01110000011,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m000111_0	),
Adb01110000100	(	adb01110000100,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m000111_0	),
Adb01110000101	(	adb01110000101,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m000111_0	),
Adb01110000110	(	adb01110000110,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m000111_0	),
Adb01110000111	(	adb01110000111,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m000111_0	),
Adb01110001000	(	adb01110001000,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m000111_0	),
Adb01110001001	(	adb01110001001,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m000111_0	),
Adb01110001010	(	adb01110001010,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m000111_0	),
Adb01110001011	(	adb01110001011,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m000111_0	),
Adb01110001100	(	adb01110001100,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m000111_0	),
Adb01110001101	(	adb01110001101,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m000111_0	),
Adb01110001110	(	adb01110001110,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m000111_0	),
Adb01110001111	(	adb01110001111,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m000111_0	),
Adb01110010000	(	adb01110010000,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m000111_0	),
Adb01110010001	(	adb01110010001,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m000111_0	),
Adb01110010010	(	adb01110010010,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m000111_0	),
Adb01110010011	(	adb01110010011,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m000111_0	),
Adb01110010100	(	adb01110010100,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m000111_0	),
Adb01110010101	(	adb01110010101,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m000111_0	),
Adb01110010110	(	adb01110010110,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m000111_0	),
Adb01110010111	(	adb01110010111,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m000111_0	),
Adb01110011000	(	adb01110011000,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m000111_0	),
Adb01110011001	(	adb01110011001,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m000111_0	),
Adb01110011010	(	adb01110011010,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m000111_0	),
Adb01110011011	(	adb01110011011,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m000111_0	),
Adb01110011100	(	adb01110011100,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m000111_0	),
Adb01110011101	(	adb01110011101,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m000111_0	),
Adb01110011110	(	adb01110011110,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m000111_0	),
Adb01110011111	(	adb01110011111,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m000111_0	),
Adb01110100000	(	adb01110100000,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m000111_0	),
Adb01110100001	(	adb01110100001,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m000111_0	),
Adb01110100010	(	adb01110100010,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m000111_0	),
Adb01110100011	(	adb01110100011,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m000111_0	),
Adb01110100100	(	adb01110100100,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m000111_0	),
Adb01110100101	(	adb01110100101,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m000111_0	),
Adb01110100110	(	adb01110100110,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m000111_0	),
Adb01110100111	(	adb01110100111,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m000111_0	),
Adb01110101000	(	adb01110101000,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m000111_0	),
Adb01110101001	(	adb01110101001,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m000111_0	),
Adb01110101010	(	adb01110101010,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m000111_0	),
Adb01110101011	(	adb01110101011,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m000111_0	),
Adb01110101100	(	adb01110101100,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m000111_0	),
Adb01110101101	(	adb01110101101,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m000111_0	),
Adb01110101110	(	adb01110101110,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m000111_0	),
Adb01110101111	(	adb01110101111,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m000111_0	),
Adb01110110000	(	adb01110110000,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m000111_0	),
Adb01110110001	(	adb01110110001,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m000111_0	),
Adb01110110010	(	adb01110110010,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m000111_0	),
Adb01110110011	(	adb01110110011,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m000111_0	),
Adb01110110100	(	adb01110110100,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m000111_0	),
Adb01110110101	(	adb01110110101,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m000111_0	),
Adb01110110110	(	adb01110110110,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m000111_0	),
Adb01110110111	(	adb01110110111,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m000111_0	),
Adb01110111000	(	adb01110111000,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m000111_0	),
Adb01110111001	(	adb01110111001,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m000111_0	),
Adb01110111010	(	adb01110111010,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m000111_0	),
Adb01110111011	(	adb01110111011,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m000111_0	),
Adb01110111100	(	adb01110111100,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m000111_0	),
Adb01110111101	(	adb01110111101,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m000111_0	),
Adb01110111110	(	adb01110111110,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m000111_0	),
Adb01110111111	(	adb01110111111,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m000111_0	),
Adb01111000000	(	adb01111000000,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m000111_0	),
Adb01111000001	(	adb01111000001,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m000111_0	),
Adb01111000010	(	adb01111000010,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m000111_0	),
Adb01111000011	(	adb01111000011,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m000111_0	),
Adb01111000100	(	adb01111000100,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m000111_0	),
Adb01111000101	(	adb01111000101,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m000111_0	),
Adb01111000110	(	adb01111000110,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m000111_0	),
Adb01111000111	(	adb01111000111,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m000111_0	),
Adb01111001000	(	adb01111001000,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m000111_0	),
Adb01111001001	(	adb01111001001,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m000111_0	),
Adb01111001010	(	adb01111001010,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m000111_0	),
Adb01111001011	(	adb01111001011,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m000111_0	),
Adb01111001100	(	adb01111001100,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m000111_0	),
Adb01111001101	(	adb01111001101,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m000111_0	),
Adb01111001110	(	adb01111001110,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m000111_0	),
Adb01111001111	(	adb01111001111,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m000111_0	),
Adb01111010000	(	adb01111010000,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m000111_0	),
Adb01111010001	(	adb01111010001,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m000111_0	),
Adb01111010010	(	adb01111010010,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m000111_0	),
Adb01111010011	(	adb01111010011,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m000111_0	),
Adb01111010100	(	adb01111010100,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m000111_0	),
Adb01111010101	(	adb01111010101,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m000111_0	),
Adb01111010110	(	adb01111010110,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m000111_0	),
Adb01111010111	(	adb01111010111,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m000111_0	),
Adb01111011000	(	adb01111011000,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m000111_0	),
Adb01111011001	(	adb01111011001,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m000111_0	),
Adb01111011010	(	adb01111011010,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m000111_0	),
Adb01111011011	(	adb01111011011,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m000111_0	),
Adb01111011100	(	adb01111011100,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m000111_0	),
Adb01111011101	(	adb01111011101,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m000111_0	),
Adb01111011110	(	adb01111011110,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m000111_0	),
Adb01111011111	(	adb01111011111,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m000111_0	),
Adb01111100000	(	adb01111100000,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m000111_0	),
Adb01111100001	(	adb01111100001,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m000111_0	),
Adb01111100010	(	adb01111100010,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m000111_0	),
Adb01111100011	(	adb01111100011,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m000111_0	),
Adb01111100100	(	adb01111100100,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m000111_0	),
Adb01111100101	(	adb01111100101,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m000111_0	),
Adb01111100110	(	adb01111100110,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m000111_0	),
Adb01111100111	(	adb01111100111,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m000111_0	),
Adb01111101000	(	adb01111101000,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m000111_0	),
Adb01111101001	(	adb01111101001,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m000111_0	),
Adb01111101010	(	adb01111101010,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m000111_0	),
Adb01111101011	(	adb01111101011,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m000111_0	),
Adb01111101100	(	adb01111101100,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m000111_0	),
Adb01111101101	(	adb01111101101,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m000111_0	),
Adb01111101110	(	adb01111101110,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m000111_0	),
Adb01111101111	(	adb01111101111,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m000111_0	),
Adb01111110000	(	adb01111110000,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m000111_0	),
Adb01111110001	(	adb01111110001,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m000111_0	),
Adb01111110010	(	adb01111110010,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m000111_0	),
Adb01111110011	(	adb01111110011,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m000111_0	),
Adb01111110100	(	adb01111110100,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m000111_0	),
Adb01111110101	(	adb01111110101,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m000111_0	),
Adb01111110110	(	adb01111110110,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m000111_0	),
Adb01111110111	(	adb01111110111,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m000111_0	),
Adb01111111000	(	adb01111111000,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m000111_0	),
Adb01111111001	(	adb01111111001,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m000111_0	),
Adb01111111010	(	adb01111111010,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m000111_0	),
Adb01111111011	(	adb01111111011,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m000111_0	),
Adb01111111100	(	adb01111111100,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m000111_0	),
Adb01111111101	(	adb01111111101,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m000111_0	),
Adb01111111110	(	adb01111111110,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m000111_0	),
Adb01111111111	(	adb01111111111,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m000111_0	),
       Adb100(adb100,n0011,n0010,n0009,dbv1),
       Adb101(adb101,n0011,n0010,m0009,dbv0),
       Adb110(adb110,n0011,m0010,n0009,m0018),
       Adb111(adb111,n0011,m0010,m0009,dbv0),
Adb10000000000	(	adb10000000000,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m111110_0	),
Adb10000000001	(	adb10000000001,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m111110_0	),
Adb10000000010	(	adb10000000010,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m111110_0	),
Adb10000000011	(	adb10000000011,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m111110_0	),
Adb10000000100	(	adb10000000100,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m111110_0	),
Adb10000000101	(	adb10000000101,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m111110_0	),
Adb10000000110	(	adb10000000110,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m111110_0	),
Adb10000000111	(	adb10000000111,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m111110_0	),
Adb10000001000	(	adb10000001000,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m111110_0	),
Adb10000001001	(	adb10000001001,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m111110_0	),
Adb10000001010	(	adb10000001010,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m111110_0	),
Adb10000001011	(	adb10000001011,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m111110_0	),
Adb10000001100	(	adb10000001100,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m111110_0	),
Adb10000001101	(	adb10000001101,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m111110_0	),
Adb10000001110	(	adb10000001110,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m111110_0	),
Adb10000001111	(	adb10000001111,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m111110_0	),
Adb10000010000	(	adb10000010000,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m111110_0	),
Adb10000010001	(	adb10000010001,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m111110_0	),
Adb10000010010	(	adb10000010010,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m111110_0	),
Adb10000010011	(	adb10000010011,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m111110_0	),
Adb10000010100	(	adb10000010100,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m111110_0	),
Adb10000010101	(	adb10000010101,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m111110_0	),
Adb10000010110	(	adb10000010110,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m111110_0	),
Adb10000010111	(	adb10000010111,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m111110_0	),
Adb10000011000	(	adb10000011000,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m111110_0	),
Adb10000011001	(	adb10000011001,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m111110_0	),
Adb10000011010	(	adb10000011010,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m111110_0	),
Adb10000011011	(	adb10000011011,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m111110_0	),
Adb10000011100	(	adb10000011100,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m111110_0	),
Adb10000011101	(	adb10000011101,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m111110_0	),
Adb10000011110	(	adb10000011110,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m111110_0	),
Adb10000011111	(	adb10000011111,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m111110_0	),
Adb10000100000	(	adb10000100000,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m111110_0	),
Adb10000100001	(	adb10000100001,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m111110_0	),
Adb10000100010	(	adb10000100010,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m111110_0	),
Adb10000100011	(	adb10000100011,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m111110_0	),
Adb10000100100	(	adb10000100100,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m111110_0	),
Adb10000100101	(	adb10000100101,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m111110_0	),
Adb10000100110	(	adb10000100110,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m111110_0	),
Adb10000100111	(	adb10000100111,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m111110_0	),
Adb10000101000	(	adb10000101000,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m111110_0	),
Adb10000101001	(	adb10000101001,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m111110_0	),
Adb10000101010	(	adb10000101010,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m111110_0	),
Adb10000101011	(	adb10000101011,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m111110_0	),
Adb10000101100	(	adb10000101100,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m111110_0	),
Adb10000101101	(	adb10000101101,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m111110_0	),
Adb10000101110	(	adb10000101110,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m111110_0	),
Adb10000101111	(	adb10000101111,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m111110_0	),
Adb10000110000	(	adb10000110000,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m111110_0	),
Adb10000110001	(	adb10000110001,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m111110_0	),
Adb10000110010	(	adb10000110010,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m111110_0	),
Adb10000110011	(	adb10000110011,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m111110_0	),
Adb10000110100	(	adb10000110100,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m111110_0	),
Adb10000110101	(	adb10000110101,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m111110_0	),
Adb10000110110	(	adb10000110110,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m111110_0	),
Adb10000110111	(	adb10000110111,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m111110_0	),
Adb10000111000	(	adb10000111000,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m111110_0	),
Adb10000111001	(	adb10000111001,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m111110_0	),
Adb10000111010	(	adb10000111010,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m111110_0	),
Adb10000111011	(	adb10000111011,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m111110_0	),
Adb10000111100	(	adb10000111100,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m111110_0	),
Adb10000111101	(	adb10000111101,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m111110_0	),
Adb10000111110	(	adb10000111110,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m111110_0	),
Adb10000111111	(	adb10000111111,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m111110_0	),
Adb10001000000	(	adb10001000000,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m111110_0	),
Adb10001000001	(	adb10001000001,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m111110_0	),
Adb10001000010	(	adb10001000010,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m111110_0	),
Adb10001000011	(	adb10001000011,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m111110_0	),
Adb10001000100	(	adb10001000100,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m111110_0	),
Adb10001000101	(	adb10001000101,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m111110_0	),
Adb10001000110	(	adb10001000110,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m111110_0	),
Adb10001000111	(	adb10001000111,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m111110_0	),
Adb10001001000	(	adb10001001000,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m111110_0	),
Adb10001001001	(	adb10001001001,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m111110_0	),
Adb10001001010	(	adb10001001010,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m111110_0	),
Adb10001001011	(	adb10001001011,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m111110_0	),
Adb10001001100	(	adb10001001100,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m111110_0	),
Adb10001001101	(	adb10001001101,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m111110_0	),
Adb10001001110	(	adb10001001110,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m111110_0	),
Adb10001001111	(	adb10001001111,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m111110_0	),
Adb10001010000	(	adb10001010000,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m111110_0	),
Adb10001010001	(	adb10001010001,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m111110_0	),
Adb10001010010	(	adb10001010010,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m111110_0	),
Adb10001010011	(	adb10001010011,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m111110_0	),
Adb10001010100	(	adb10001010100,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m111110_0	),
Adb10001010101	(	adb10001010101,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m111110_0	),
Adb10001010110	(	adb10001010110,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m111110_0	),
Adb10001010111	(	adb10001010111,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m111110_0	),
Adb10001011000	(	adb10001011000,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m111110_0	),
Adb10001011001	(	adb10001011001,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m111110_0	),
Adb10001011010	(	adb10001011010,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m111110_0	),
Adb10001011011	(	adb10001011011,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m111110_0	),
Adb10001011100	(	adb10001011100,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m111110_0	),
Adb10001011101	(	adb10001011101,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m111110_0	),
Adb10001011110	(	adb10001011110,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m111110_0	),
Adb10001011111	(	adb10001011111,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m111110_0	),
Adb10001100000	(	adb10001100000,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m111110_0	),
Adb10001100001	(	adb10001100001,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m111110_0	),
Adb10001100010	(	adb10001100010,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m111110_0	),
Adb10001100011	(	adb10001100011,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m111110_0	),
Adb10001100100	(	adb10001100100,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m111110_0	),
Adb10001100101	(	adb10001100101,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m111110_0	),
Adb10001100110	(	adb10001100110,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m111110_0	),
Adb10001100111	(	adb10001100111,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m111110_0	),
Adb10001101000	(	adb10001101000,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m111110_0	),
Adb10001101001	(	adb10001101001,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m111110_0	),
Adb10001101010	(	adb10001101010,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m111110_0	),
Adb10001101011	(	adb10001101011,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m111110_0	),
Adb10001101100	(	adb10001101100,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m111110_0	),
Adb10001101101	(	adb10001101101,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m111110_0	),
Adb10001101110	(	adb10001101110,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m111110_0	),
Adb10001101111	(	adb10001101111,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m111110_0	),
Adb10001110000	(	adb10001110000,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m111110_0	),
Adb10001110001	(	adb10001110001,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m111110_0	),
Adb10001110010	(	adb10001110010,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m111110_0	),
Adb10001110011	(	adb10001110011,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m111110_0	),
Adb10001110100	(	adb10001110100,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m111110_0	),
Adb10001110101	(	adb10001110101,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m111110_0	),
Adb10001110110	(	adb10001110110,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m111110_0	),
Adb10001110111	(	adb10001110111,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m111110_0	),
Adb10001111000	(	adb10001111000,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m111110_0	),
Adb10001111001	(	adb10001111001,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m111110_0	),
Adb10001111010	(	adb10001111010,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m111110_0	),
Adb10001111011	(	adb10001111011,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m111110_0	),
Adb10001111100	(	adb10001111100,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m111110_0	),
Adb10001111101	(	adb10001111101,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m111110_0	),
Adb10001111110	(	adb10001111110,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m111110_0	),
Adb10001111111	(	adb10001111111,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m111110_0	),
Adb10010000000	(	adb10010000000,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m110110_0	),
Adb10010000001	(	adb10010000001,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m110110_0	),
Adb10010000010	(	adb10010000010,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m110110_0	),
Adb10010000011	(	adb10010000011,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m110110_0	),
Adb10010000100	(	adb10010000100,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m110110_0	),
Adb10010000101	(	adb10010000101,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m110110_0	),
Adb10010000110	(	adb10010000110,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m110110_0	),
Adb10010000111	(	adb10010000111,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m110110_0	),
Adb10010001000	(	adb10010001000,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m110110_0	),
Adb10010001001	(	adb10010001001,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m110110_0	),
Adb10010001010	(	adb10010001010,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m110110_0	),
Adb10010001011	(	adb10010001011,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m110110_0	),
Adb10010001100	(	adb10010001100,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m110110_0	),
Adb10010001101	(	adb10010001101,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m110110_0	),
Adb10010001110	(	adb10010001110,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m110110_0	),
Adb10010001111	(	adb10010001111,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m110110_0	),
Adb10010010000	(	adb10010010000,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m110110_0	),
Adb10010010001	(	adb10010010001,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m110110_0	),
Adb10010010010	(	adb10010010010,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m110110_0	),
Adb10010010011	(	adb10010010011,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m110110_0	),
Adb10010010100	(	adb10010010100,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m110110_0	),
Adb10010010101	(	adb10010010101,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m110110_0	),
Adb10010010110	(	adb10010010110,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m110110_0	),
Adb10010010111	(	adb10010010111,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m110110_0	),
Adb10010011000	(	adb10010011000,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m110110_0	),
Adb10010011001	(	adb10010011001,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m110110_0	),
Adb10010011010	(	adb10010011010,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m110110_0	),
Adb10010011011	(	adb10010011011,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m110110_0	),
Adb10010011100	(	adb10010011100,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m110110_0	),
Adb10010011101	(	adb10010011101,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m110110_0	),
Adb10010011110	(	adb10010011110,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m110110_0	),
Adb10010011111	(	adb10010011111,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m110110_0	),
Adb10010100000	(	adb10010100000,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m110110_0	),
Adb10010100001	(	adb10010100001,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m110110_0	),
Adb10010100010	(	adb10010100010,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m110110_0	),
Adb10010100011	(	adb10010100011,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m110110_0	),
Adb10010100100	(	adb10010100100,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m110110_0	),
Adb10010100101	(	adb10010100101,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m110110_0	),
Adb10010100110	(	adb10010100110,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m110110_0	),
Adb10010100111	(	adb10010100111,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m110110_0	),
Adb10010101000	(	adb10010101000,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m110110_0	),
Adb10010101001	(	adb10010101001,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m110110_0	),
Adb10010101010	(	adb10010101010,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m110110_0	),
Adb10010101011	(	adb10010101011,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m110110_0	),
Adb10010101100	(	adb10010101100,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m110110_0	),
Adb10010101101	(	adb10010101101,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m110110_0	),
Adb10010101110	(	adb10010101110,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m110110_0	),
Adb10010101111	(	adb10010101111,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m110110_0	),
Adb10010110000	(	adb10010110000,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m110110_0	),
Adb10010110001	(	adb10010110001,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m110110_0	),
Adb10010110010	(	adb10010110010,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m110110_0	),
Adb10010110011	(	adb10010110011,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m110110_0	),
Adb10010110100	(	adb10010110100,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m110110_0	),
Adb10010110101	(	adb10010110101,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m110110_0	),
Adb10010110110	(	adb10010110110,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m110110_0	),
Adb10010110111	(	adb10010110111,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m110110_0	),
Adb10010111000	(	adb10010111000,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m110110_0	),
Adb10010111001	(	adb10010111001,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m110110_0	),
Adb10010111010	(	adb10010111010,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m110110_0	),
Adb10010111011	(	adb10010111011,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m110110_0	),
Adb10010111100	(	adb10010111100,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m110110_0	),
Adb10010111101	(	adb10010111101,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m110110_0	),
Adb10010111110	(	adb10010111110,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m110110_0	),
Adb10010111111	(	adb10010111111,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m110110_0	),
Adb10011000000	(	adb10011000000,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m110110_0	),
Adb10011000001	(	adb10011000001,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m110110_0	),
Adb10011000010	(	adb10011000010,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m110110_0	),
Adb10011000011	(	adb10011000011,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m110110_0	),
Adb10011000100	(	adb10011000100,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m110110_0	),
Adb10011000101	(	adb10011000101,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m110110_0	),
Adb10011000110	(	adb10011000110,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m110110_0	),
Adb10011000111	(	adb10011000111,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m110110_0	),
Adb10011001000	(	adb10011001000,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m110110_0	),
Adb10011001001	(	adb10011001001,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m110110_0	),
Adb10011001010	(	adb10011001010,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m110110_0	),
Adb10011001011	(	adb10011001011,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m110110_0	),
Adb10011001100	(	adb10011001100,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m110110_0	),
Adb10011001101	(	adb10011001101,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m110110_0	),
Adb10011001110	(	adb10011001110,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m110110_0	),
Adb10011001111	(	adb10011001111,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m110110_0	),
Adb10011010000	(	adb10011010000,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m110110_0	),
Adb10011010001	(	adb10011010001,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m110110_0	),
Adb10011010010	(	adb10011010010,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m110110_0	),
Adb10011010011	(	adb10011010011,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m110110_0	),
Adb10011010100	(	adb10011010100,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m110110_0	),
Adb10011010101	(	adb10011010101,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m110110_0	),
Adb10011010110	(	adb10011010110,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m110110_0	),
Adb10011010111	(	adb10011010111,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m110110_0	),
Adb10011011000	(	adb10011011000,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m110110_0	),
Adb10011011001	(	adb10011011001,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m110110_0	),
Adb10011011010	(	adb10011011010,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m110110_0	),
Adb10011011011	(	adb10011011011,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m110110_0	),
Adb10011011100	(	adb10011011100,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m110110_0	),
Adb10011011101	(	adb10011011101,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m110110_0	),
Adb10011011110	(	adb10011011110,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m110110_0	),
Adb10011011111	(	adb10011011111,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m110110_0	),
Adb10011100000	(	adb10011100000,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m110110_0	),
Adb10011100001	(	adb10011100001,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m110110_0	),
Adb10011100010	(	adb10011100010,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m110110_0	),
Adb10011100011	(	adb10011100011,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m110110_0	),
Adb10011100100	(	adb10011100100,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m110110_0	),
Adb10011100101	(	adb10011100101,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m110110_0	),
Adb10011100110	(	adb10011100110,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m110110_0	),
Adb10011100111	(	adb10011100111,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m110110_0	),
Adb10011101000	(	adb10011101000,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m110110_0	),
Adb10011101001	(	adb10011101001,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m110110_0	),
Adb10011101010	(	adb10011101010,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m110110_0	),
Adb10011101011	(	adb10011101011,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m110110_0	),
Adb10011101100	(	adb10011101100,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m110110_0	),
Adb10011101101	(	adb10011101101,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m110110_0	),
Adb10011101110	(	adb10011101110,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m110110_0	),
Adb10011101111	(	adb10011101111,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m110110_0	),
Adb10011110000	(	adb10011110000,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m110110_0	),
Adb10011110001	(	adb10011110001,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m110110_0	),
Adb10011110010	(	adb10011110010,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m110110_0	),
Adb10011110011	(	adb10011110011,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m110110_0	),
Adb10011110100	(	adb10011110100,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m110110_0	),
Adb10011110101	(	adb10011110101,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m110110_0	),
Adb10011110110	(	adb10011110110,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m110110_0	),
Adb10011110111	(	adb10011110111,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m110110_0	),
Adb10011111000	(	adb10011111000,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m110110_0	),
Adb10011111001	(	adb10011111001,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m110110_0	),
Adb10011111010	(	adb10011111010,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m110110_0	),
Adb10011111011	(	adb10011111011,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m110110_0	),
Adb10011111100	(	adb10011111100,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m110110_0	),
Adb10011111101	(	adb10011111101,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m110110_0	),
Adb10011111110	(	adb10011111110,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m110110_0	),
Adb10011111111	(	adb10011111111,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m110110_0	),
Adb10100000000	(	adb10100000000,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m101110_0	),
Adb10100000001	(	adb10100000001,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m101110_0	),
Adb10100000010	(	adb10100000010,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m101110_0	),
Adb10100000011	(	adb10100000011,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m101110_0	),
Adb10100000100	(	adb10100000100,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m101110_0	),
Adb10100000101	(	adb10100000101,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m101110_0	),
Adb10100000110	(	adb10100000110,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m101110_0	),
Adb10100000111	(	adb10100000111,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m101110_0	),
Adb10100001000	(	adb10100001000,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m101110_0	),
Adb10100001001	(	adb10100001001,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m101110_0	),
Adb10100001010	(	adb10100001010,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m101110_0	),
Adb10100001011	(	adb10100001011,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m101110_0	),
Adb10100001100	(	adb10100001100,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m101110_0	),
Adb10100001101	(	adb10100001101,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m101110_0	),
Adb10100001110	(	adb10100001110,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m101110_0	),
Adb10100001111	(	adb10100001111,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m101110_0	),
Adb10100010000	(	adb10100010000,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m101110_0	),
Adb10100010001	(	adb10100010001,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m101110_0	),
Adb10100010010	(	adb10100010010,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m101110_0	),
Adb10100010011	(	adb10100010011,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m101110_0	),
Adb10100010100	(	adb10100010100,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m101110_0	),
Adb10100010101	(	adb10100010101,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m101110_0	),
Adb10100010110	(	adb10100010110,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m101110_0	),
Adb10100010111	(	adb10100010111,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m101110_0	),
Adb10100011000	(	adb10100011000,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m101110_0	),
Adb10100011001	(	adb10100011001,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m101110_0	),
Adb10100011010	(	adb10100011010,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m101110_0	),
Adb10100011011	(	adb10100011011,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m101110_0	),
Adb10100011100	(	adb10100011100,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m101110_0	),
Adb10100011101	(	adb10100011101,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m101110_0	),
Adb10100011110	(	adb10100011110,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m101110_0	),
Adb10100011111	(	adb10100011111,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m101110_0	),
Adb10100100000	(	adb10100100000,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m101110_0	),
Adb10100100001	(	adb10100100001,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m101110_0	),
Adb10100100010	(	adb10100100010,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m101110_0	),
Adb10100100011	(	adb10100100011,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m101110_0	),
Adb10100100100	(	adb10100100100,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m101110_0	),
Adb10100100101	(	adb10100100101,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m101110_0	),
Adb10100100110	(	adb10100100110,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m101110_0	),
Adb10100100111	(	adb10100100111,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m101110_0	),
Adb10100101000	(	adb10100101000,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m101110_0	),
Adb10100101001	(	adb10100101001,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m101110_0	),
Adb10100101010	(	adb10100101010,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m101110_0	),
Adb10100101011	(	adb10100101011,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m101110_0	),
Adb10100101100	(	adb10100101100,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m101110_0	),
Adb10100101101	(	adb10100101101,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m101110_0	),
Adb10100101110	(	adb10100101110,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m101110_0	),
Adb10100101111	(	adb10100101111,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m101110_0	),
Adb10100110000	(	adb10100110000,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m101110_0	),
Adb10100110001	(	adb10100110001,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m101110_0	),
Adb10100110010	(	adb10100110010,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m101110_0	),
Adb10100110011	(	adb10100110011,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m101110_0	),
Adb10100110100	(	adb10100110100,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m101110_0	),
Adb10100110101	(	adb10100110101,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m101110_0	),
Adb10100110110	(	adb10100110110,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m101110_0	),
Adb10100110111	(	adb10100110111,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m101110_0	),
Adb10100111000	(	adb10100111000,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m101110_0	),
Adb10100111001	(	adb10100111001,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m101110_0	),
Adb10100111010	(	adb10100111010,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m101110_0	),
Adb10100111011	(	adb10100111011,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m101110_0	),
Adb10100111100	(	adb10100111100,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m101110_0	),
Adb10100111101	(	adb10100111101,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m101110_0	),
Adb10100111110	(	adb10100111110,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m101110_0	),
Adb10100111111	(	adb10100111111,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m101110_0	),
Adb10101000000	(	adb10101000000,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m101110_0	),
Adb10101000001	(	adb10101000001,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m101110_0	),
Adb10101000010	(	adb10101000010,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m101110_0	),
Adb10101000011	(	adb10101000011,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m101110_0	),
Adb10101000100	(	adb10101000100,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m101110_0	),
Adb10101000101	(	adb10101000101,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m101110_0	),
Adb10101000110	(	adb10101000110,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m101110_0	),
Adb10101000111	(	adb10101000111,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m101110_0	),
Adb10101001000	(	adb10101001000,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m101110_0	),
Adb10101001001	(	adb10101001001,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m101110_0	),
Adb10101001010	(	adb10101001010,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m101110_0	),
Adb10101001011	(	adb10101001011,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m101110_0	),
Adb10101001100	(	adb10101001100,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m101110_0	),
Adb10101001101	(	adb10101001101,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m101110_0	),
Adb10101001110	(	adb10101001110,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m101110_0	),
Adb10101001111	(	adb10101001111,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m101110_0	),
Adb10101010000	(	adb10101010000,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m101110_0	),
Adb10101010001	(	adb10101010001,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m101110_0	),
Adb10101010010	(	adb10101010010,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m101110_0	),
Adb10101010011	(	adb10101010011,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m101110_0	),
Adb10101010100	(	adb10101010100,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m101110_0	),
Adb10101010101	(	adb10101010101,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m101110_0	),
Adb10101010110	(	adb10101010110,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m101110_0	),
Adb10101010111	(	adb10101010111,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m101110_0	),
Adb10101011000	(	adb10101011000,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m101110_0	),
Adb10101011001	(	adb10101011001,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m101110_0	),
Adb10101011010	(	adb10101011010,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m101110_0	),
Adb10101011011	(	adb10101011011,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m101110_0	),
Adb10101011100	(	adb10101011100,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m101110_0	),
Adb10101011101	(	adb10101011101,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m101110_0	),
Adb10101011110	(	adb10101011110,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m101110_0	),
Adb10101011111	(	adb10101011111,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m101110_0	),
Adb10101100000	(	adb10101100000,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m101110_0	),
Adb10101100001	(	adb10101100001,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m101110_0	),
Adb10101100010	(	adb10101100010,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m101110_0	),
Adb10101100011	(	adb10101100011,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m101110_0	),
Adb10101100100	(	adb10101100100,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m101110_0	),
Adb10101100101	(	adb10101100101,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m101110_0	),
Adb10101100110	(	adb10101100110,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m101110_0	),
Adb10101100111	(	adb10101100111,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m101110_0	),
Adb10101101000	(	adb10101101000,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m101110_0	),
Adb10101101001	(	adb10101101001,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m101110_0	),
Adb10101101010	(	adb10101101010,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m101110_0	),
Adb10101101011	(	adb10101101011,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m101110_0	),
Adb10101101100	(	adb10101101100,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m101110_0	),
Adb10101101101	(	adb10101101101,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m101110_0	),
Adb10101101110	(	adb10101101110,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m101110_0	),
Adb10101101111	(	adb10101101111,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m101110_0	),
Adb10101110000	(	adb10101110000,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m101110_0	),
Adb10101110001	(	adb10101110001,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m101110_0	),
Adb10101110010	(	adb10101110010,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m101110_0	),
Adb10101110011	(	adb10101110011,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m101110_0	),
Adb10101110100	(	adb10101110100,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m101110_0	),
Adb10101110101	(	adb10101110101,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m101110_0	),
Adb10101110110	(	adb10101110110,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m101110_0	),
Adb10101110111	(	adb10101110111,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m101110_0	),
Adb10101111000	(	adb10101111000,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m101110_0	),
Adb10101111001	(	adb10101111001,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m101110_0	),
Adb10101111010	(	adb10101111010,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m101110_0	),
Adb10101111011	(	adb10101111011,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m101110_0	),
Adb10101111100	(	adb10101111100,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m101110_0	),
Adb10101111101	(	adb10101111101,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m101110_0	),
Adb10101111110	(	adb10101111110,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m101110_0	),
Adb10101111111	(	adb10101111111,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m101110_0	),
Adb10110000000	(	adb10110000000,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m100110_0	),
Adb10110000001	(	adb10110000001,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m100110_0	),
Adb10110000010	(	adb10110000010,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m100110_0	),
Adb10110000011	(	adb10110000011,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m100110_0	),
Adb10110000100	(	adb10110000100,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m100110_0	),
Adb10110000101	(	adb10110000101,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m100110_0	),
Adb10110000110	(	adb10110000110,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m100110_0	),
Adb10110000111	(	adb10110000111,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m100110_0	),
Adb10110001000	(	adb10110001000,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m100110_0	),
Adb10110001001	(	adb10110001001,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m100110_0	),
Adb10110001010	(	adb10110001010,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m100110_0	),
Adb10110001011	(	adb10110001011,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m100110_0	),
Adb10110001100	(	adb10110001100,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m100110_0	),
Adb10110001101	(	adb10110001101,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m100110_0	),
Adb10110001110	(	adb10110001110,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m100110_0	),
Adb10110001111	(	adb10110001111,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m100110_0	),
Adb10110010000	(	adb10110010000,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m100110_0	),
Adb10110010001	(	adb10110010001,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m100110_0	),
Adb10110010010	(	adb10110010010,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m100110_0	),
Adb10110010011	(	adb10110010011,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m100110_0	),
Adb10110010100	(	adb10110010100,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m100110_0	),
Adb10110010101	(	adb10110010101,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m100110_0	),
Adb10110010110	(	adb10110010110,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m100110_0	),
Adb10110010111	(	adb10110010111,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m100110_0	),
Adb10110011000	(	adb10110011000,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m100110_0	),
Adb10110011001	(	adb10110011001,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m100110_0	),
Adb10110011010	(	adb10110011010,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m100110_0	),
Adb10110011011	(	adb10110011011,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m100110_0	),
Adb10110011100	(	adb10110011100,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m100110_0	),
Adb10110011101	(	adb10110011101,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m100110_0	),
Adb10110011110	(	adb10110011110,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m100110_0	),
Adb10110011111	(	adb10110011111,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m100110_0	),
Adb10110100000	(	adb10110100000,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m100110_0	),
Adb10110100001	(	adb10110100001,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m100110_0	),
Adb10110100010	(	adb10110100010,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m100110_0	),
Adb10110100011	(	adb10110100011,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m100110_0	),
Adb10110100100	(	adb10110100100,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m100110_0	),
Adb10110100101	(	adb10110100101,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m100110_0	),
Adb10110100110	(	adb10110100110,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m100110_0	),
Adb10110100111	(	adb10110100111,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m100110_0	),
Adb10110101000	(	adb10110101000,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m100110_0	),
Adb10110101001	(	adb10110101001,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m100110_0	),
Adb10110101010	(	adb10110101010,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m100110_0	),
Adb10110101011	(	adb10110101011,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m100110_0	),
Adb10110101100	(	adb10110101100,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m100110_0	),
Adb10110101101	(	adb10110101101,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m100110_0	),
Adb10110101110	(	adb10110101110,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m100110_0	),
Adb10110101111	(	adb10110101111,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m100110_0	),
Adb10110110000	(	adb10110110000,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m100110_0	),
Adb10110110001	(	adb10110110001,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m100110_0	),
Adb10110110010	(	adb10110110010,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m100110_0	),
Adb10110110011	(	adb10110110011,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m100110_0	),
Adb10110110100	(	adb10110110100,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m100110_0	),
Adb10110110101	(	adb10110110101,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m100110_0	),
Adb10110110110	(	adb10110110110,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m100110_0	),
Adb10110110111	(	adb10110110111,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m100110_0	),
Adb10110111000	(	adb10110111000,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m100110_0	),
Adb10110111001	(	adb10110111001,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m100110_0	),
Adb10110111010	(	adb10110111010,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m100110_0	),
Adb10110111011	(	adb10110111011,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m100110_0	),
Adb10110111100	(	adb10110111100,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m100110_0	),
Adb10110111101	(	adb10110111101,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m100110_0	),
Adb10110111110	(	adb10110111110,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m100110_0	),
Adb10110111111	(	adb10110111111,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m100110_0	),
Adb10111000000	(	adb10111000000,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m100110_0	),
Adb10111000001	(	adb10111000001,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m100110_0	),
Adb10111000010	(	adb10111000010,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m100110_0	),
Adb10111000011	(	adb10111000011,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m100110_0	),
Adb10111000100	(	adb10111000100,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m100110_0	),
Adb10111000101	(	adb10111000101,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m100110_0	),
Adb10111000110	(	adb10111000110,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m100110_0	),
Adb10111000111	(	adb10111000111,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m100110_0	),
Adb10111001000	(	adb10111001000,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m100110_0	),
Adb10111001001	(	adb10111001001,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m100110_0	),
Adb10111001010	(	adb10111001010,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m100110_0	),
Adb10111001011	(	adb10111001011,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m100110_0	),
Adb10111001100	(	adb10111001100,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m100110_0	),
Adb10111001101	(	adb10111001101,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m100110_0	),
Adb10111001110	(	adb10111001110,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m100110_0	),
Adb10111001111	(	adb10111001111,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m100110_0	),
Adb10111010000	(	adb10111010000,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m100110_0	),
Adb10111010001	(	adb10111010001,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m100110_0	),
Adb10111010010	(	adb10111010010,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m100110_0	),
Adb10111010011	(	adb10111010011,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m100110_0	),
Adb10111010100	(	adb10111010100,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m100110_0	),
Adb10111010101	(	adb10111010101,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m100110_0	),
Adb10111010110	(	adb10111010110,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m100110_0	),
Adb10111010111	(	adb10111010111,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m100110_0	),
Adb10111011000	(	adb10111011000,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m100110_0	),
Adb10111011001	(	adb10111011001,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m100110_0	),
Adb10111011010	(	adb10111011010,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m100110_0	),
Adb10111011011	(	adb10111011011,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m100110_0	),
Adb10111011100	(	adb10111011100,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m100110_0	),
Adb10111011101	(	adb10111011101,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m100110_0	),
Adb10111011110	(	adb10111011110,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m100110_0	),
Adb10111011111	(	adb10111011111,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m100110_0	),
Adb10111100000	(	adb10111100000,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m100110_0	),
Adb10111100001	(	adb10111100001,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m100110_0	),
Adb10111100010	(	adb10111100010,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m100110_0	),
Adb10111100011	(	adb10111100011,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m100110_0	),
Adb10111100100	(	adb10111100100,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m100110_0	),
Adb10111100101	(	adb10111100101,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m100110_0	),
Adb10111100110	(	adb10111100110,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m100110_0	),
Adb10111100111	(	adb10111100111,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m100110_0	),
Adb10111101000	(	adb10111101000,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m100110_0	),
Adb10111101001	(	adb10111101001,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m100110_0	),
Adb10111101010	(	adb10111101010,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m100110_0	),
Adb10111101011	(	adb10111101011,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m100110_0	),
Adb10111101100	(	adb10111101100,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m100110_0	),
Adb10111101101	(	adb10111101101,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m100110_0	),
Adb10111101110	(	adb10111101110,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m100110_0	),
Adb10111101111	(	adb10111101111,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m100110_0	),
Adb10111110000	(	adb10111110000,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m100110_0	),
Adb10111110001	(	adb10111110001,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m100110_0	),
Adb10111110010	(	adb10111110010,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m100110_0	),
Adb10111110011	(	adb10111110011,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m100110_0	),
Adb10111110100	(	adb10111110100,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m100110_0	),
Adb10111110101	(	adb10111110101,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m100110_0	),
Adb10111110110	(	adb10111110110,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m100110_0	),
Adb10111110111	(	adb10111110111,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m100110_0	),
Adb10111111000	(	adb10111111000,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m100110_0	),
Adb10111111001	(	adb10111111001,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m100110_0	),
Adb10111111010	(	adb10111111010,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m100110_0	),
Adb10111111011	(	adb10111111011,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m100110_0	),
Adb10111111100	(	adb10111111100,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m100110_0	),
Adb10111111101	(	adb10111111101,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m100110_0	),
Adb10111111110	(	adb10111111110,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m100110_0	),
Adb10111111111	(	adb10111111111,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m100110_0	),
Adb11000000000	(	adb11000000000,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m011110_0	),
Adb11000000001	(	adb11000000001,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m011110_0	),
Adb11000000010	(	adb11000000010,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m011110_0	),
Adb11000000011	(	adb11000000011,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m011110_0	),
Adb11000000100	(	adb11000000100,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m011110_0	),
Adb11000000101	(	adb11000000101,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m011110_0	),
Adb11000000110	(	adb11000000110,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m011110_0	),
Adb11000000111	(	adb11000000111,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m011110_0	),
Adb11000001000	(	adb11000001000,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m011110_0	),
Adb11000001001	(	adb11000001001,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m011110_0	),
Adb11000001010	(	adb11000001010,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m011110_0	),
Adb11000001011	(	adb11000001011,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m011110_0	),
Adb11000001100	(	adb11000001100,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m011110_0	),
Adb11000001101	(	adb11000001101,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m011110_0	),
Adb11000001110	(	adb11000001110,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m011110_0	),
Adb11000001111	(	adb11000001111,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m011110_0	),
Adb11000010000	(	adb11000010000,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m011110_0	),
Adb11000010001	(	adb11000010001,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m011110_0	),
Adb11000010010	(	adb11000010010,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m011110_0	),
Adb11000010011	(	adb11000010011,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m011110_0	),
Adb11000010100	(	adb11000010100,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m011110_0	),
Adb11000010101	(	adb11000010101,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m011110_0	),
Adb11000010110	(	adb11000010110,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m011110_0	),
Adb11000010111	(	adb11000010111,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m011110_0	),
Adb11000011000	(	adb11000011000,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m011110_0	),
Adb11000011001	(	adb11000011001,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m011110_0	),
Adb11000011010	(	adb11000011010,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m011110_0	),
Adb11000011011	(	adb11000011011,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m011110_0	),
Adb11000011100	(	adb11000011100,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m011110_0	),
Adb11000011101	(	adb11000011101,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m011110_0	),
Adb11000011110	(	adb11000011110,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m011110_0	),
Adb11000011111	(	adb11000011111,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m011110_0	),
Adb11000100000	(	adb11000100000,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m011110_0	),
Adb11000100001	(	adb11000100001,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m011110_0	),
Adb11000100010	(	adb11000100010,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m011110_0	),
Adb11000100011	(	adb11000100011,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m011110_0	),
Adb11000100100	(	adb11000100100,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m011110_0	),
Adb11000100101	(	adb11000100101,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m011110_0	),
Adb11000100110	(	adb11000100110,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m011110_0	),
Adb11000100111	(	adb11000100111,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m011110_0	),
Adb11000101000	(	adb11000101000,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m011110_0	),
Adb11000101001	(	adb11000101001,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m011110_0	),
Adb11000101010	(	adb11000101010,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m011110_0	),
Adb11000101011	(	adb11000101011,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m011110_0	),
Adb11000101100	(	adb11000101100,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m011110_0	),
Adb11000101101	(	adb11000101101,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m011110_0	),
Adb11000101110	(	adb11000101110,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m011110_0	),
Adb11000101111	(	adb11000101111,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m011110_0	),
Adb11000110000	(	adb11000110000,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m011110_0	),
Adb11000110001	(	adb11000110001,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m011110_0	),
Adb11000110010	(	adb11000110010,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m011110_0	),
Adb11000110011	(	adb11000110011,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m011110_0	),
Adb11000110100	(	adb11000110100,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m011110_0	),
Adb11000110101	(	adb11000110101,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m011110_0	),
Adb11000110110	(	adb11000110110,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m011110_0	),
Adb11000110111	(	adb11000110111,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m011110_0	),
Adb11000111000	(	adb11000111000,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m011110_0	),
Adb11000111001	(	adb11000111001,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m011110_0	),
Adb11000111010	(	adb11000111010,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m011110_0	),
Adb11000111011	(	adb11000111011,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m011110_0	),
Adb11000111100	(	adb11000111100,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m011110_0	),
Adb11000111101	(	adb11000111101,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m011110_0	),
Adb11000111110	(	adb11000111110,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m011110_0	),
Adb11000111111	(	adb11000111111,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m011110_0	),
Adb11001000000	(	adb11001000000,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m011110_0	),
Adb11001000001	(	adb11001000001,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m011110_0	),
Adb11001000010	(	adb11001000010,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m011110_0	),
Adb11001000011	(	adb11001000011,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m011110_0	),
Adb11001000100	(	adb11001000100,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m011110_0	),
Adb11001000101	(	adb11001000101,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m011110_0	),
Adb11001000110	(	adb11001000110,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m011110_0	),
Adb11001000111	(	adb11001000111,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m011110_0	),
Adb11001001000	(	adb11001001000,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m011110_0	),
Adb11001001001	(	adb11001001001,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m011110_0	),
Adb11001001010	(	adb11001001010,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m011110_0	),
Adb11001001011	(	adb11001001011,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m011110_0	),
Adb11001001100	(	adb11001001100,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m011110_0	),
Adb11001001101	(	adb11001001101,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m011110_0	),
Adb11001001110	(	adb11001001110,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m011110_0	),
Adb11001001111	(	adb11001001111,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m011110_0	),
Adb11001010000	(	adb11001010000,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m011110_0	),
Adb11001010001	(	adb11001010001,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m011110_0	),
Adb11001010010	(	adb11001010010,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m011110_0	),
Adb11001010011	(	adb11001010011,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m011110_0	),
Adb11001010100	(	adb11001010100,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m011110_0	),
Adb11001010101	(	adb11001010101,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m011110_0	),
Adb11001010110	(	adb11001010110,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m011110_0	),
Adb11001010111	(	adb11001010111,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m011110_0	),
Adb11001011000	(	adb11001011000,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m011110_0	),
Adb11001011001	(	adb11001011001,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m011110_0	),
Adb11001011010	(	adb11001011010,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m011110_0	),
Adb11001011011	(	adb11001011011,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m011110_0	),
Adb11001011100	(	adb11001011100,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m011110_0	),
Adb11001011101	(	adb11001011101,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m011110_0	),
Adb11001011110	(	adb11001011110,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m011110_0	),
Adb11001011111	(	adb11001011111,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m011110_0	),
Adb11001100000	(	adb11001100000,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m011110_0	),
Adb11001100001	(	adb11001100001,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m011110_0	),
Adb11001100010	(	adb11001100010,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m011110_0	),
Adb11001100011	(	adb11001100011,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m011110_0	),
Adb11001100100	(	adb11001100100,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m011110_0	),
Adb11001100101	(	adb11001100101,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m011110_0	),
Adb11001100110	(	adb11001100110,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m011110_0	),
Adb11001100111	(	adb11001100111,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m011110_0	),
Adb11001101000	(	adb11001101000,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m011110_0	),
Adb11001101001	(	adb11001101001,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m011110_0	),
Adb11001101010	(	adb11001101010,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m011110_0	),
Adb11001101011	(	adb11001101011,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m011110_0	),
Adb11001101100	(	adb11001101100,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m011110_0	),
Adb11001101101	(	adb11001101101,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m011110_0	),
Adb11001101110	(	adb11001101110,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m011110_0	),
Adb11001101111	(	adb11001101111,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m011110_0	),
Adb11001110000	(	adb11001110000,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m011110_0	),
Adb11001110001	(	adb11001110001,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m011110_0	),
Adb11001110010	(	adb11001110010,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m011110_0	),
Adb11001110011	(	adb11001110011,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m011110_0	),
Adb11001110100	(	adb11001110100,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m011110_0	),
Adb11001110101	(	adb11001110101,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m011110_0	),
Adb11001110110	(	adb11001110110,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m011110_0	),
Adb11001110111	(	adb11001110111,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m011110_0	),
Adb11001111000	(	adb11001111000,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m011110_0	),
Adb11001111001	(	adb11001111001,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m011110_0	),
Adb11001111010	(	adb11001111010,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m011110_0	),
Adb11001111011	(	adb11001111011,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m011110_0	),
Adb11001111100	(	adb11001111100,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m011110_0	),
Adb11001111101	(	adb11001111101,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m011110_0	),
Adb11001111110	(	adb11001111110,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m011110_0	),
Adb11001111111	(	adb11001111111,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m011110_0	),
Adb11010000000	(	adb11010000000,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m010110_0	),
Adb11010000001	(	adb11010000001,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m010110_0	),
Adb11010000010	(	adb11010000010,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m010110_0	),
Adb11010000011	(	adb11010000011,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m010110_0	),
Adb11010000100	(	adb11010000100,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m010110_0	),
Adb11010000101	(	adb11010000101,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m010110_0	),
Adb11010000110	(	adb11010000110,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m010110_0	),
Adb11010000111	(	adb11010000111,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m010110_0	),
Adb11010001000	(	adb11010001000,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m010110_0	),
Adb11010001001	(	adb11010001001,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m010110_0	),
Adb11010001010	(	adb11010001010,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m010110_0	),
Adb11010001011	(	adb11010001011,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m010110_0	),
Adb11010001100	(	adb11010001100,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m010110_0	),
Adb11010001101	(	adb11010001101,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m010110_0	),
Adb11010001110	(	adb11010001110,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m010110_0	),
Adb11010001111	(	adb11010001111,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m010110_0	),
Adb11010010000	(	adb11010010000,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m010110_0	),
Adb11010010001	(	adb11010010001,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m010110_0	),
Adb11010010010	(	adb11010010010,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m010110_0	),
Adb11010010011	(	adb11010010011,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m010110_0	),
Adb11010010100	(	adb11010010100,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m010110_0	),
Adb11010010101	(	adb11010010101,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m010110_0	),
Adb11010010110	(	adb11010010110,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m010110_0	),
Adb11010010111	(	adb11010010111,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m010110_0	),
Adb11010011000	(	adb11010011000,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m010110_0	),
Adb11010011001	(	adb11010011001,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m010110_0	),
Adb11010011010	(	adb11010011010,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m010110_0	),
Adb11010011011	(	adb11010011011,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m010110_0	),
Adb11010011100	(	adb11010011100,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m010110_0	),
Adb11010011101	(	adb11010011101,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m010110_0	),
Adb11010011110	(	adb11010011110,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m010110_0	),
Adb11010011111	(	adb11010011111,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m010110_0	),
Adb11010100000	(	adb11010100000,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m010110_0	),
Adb11010100001	(	adb11010100001,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m010110_0	),
Adb11010100010	(	adb11010100010,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m010110_0	),
Adb11010100011	(	adb11010100011,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m010110_0	),
Adb11010100100	(	adb11010100100,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m010110_0	),
Adb11010100101	(	adb11010100101,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m010110_0	),
Adb11010100110	(	adb11010100110,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m010110_0	),
Adb11010100111	(	adb11010100111,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m010110_0	),
Adb11010101000	(	adb11010101000,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m010110_0	),
Adb11010101001	(	adb11010101001,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m010110_0	),
Adb11010101010	(	adb11010101010,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m010110_0	),
Adb11010101011	(	adb11010101011,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m010110_0	),
Adb11010101100	(	adb11010101100,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m010110_0	),
Adb11010101101	(	adb11010101101,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m010110_0	),
Adb11010101110	(	adb11010101110,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m010110_0	),
Adb11010101111	(	adb11010101111,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m010110_0	),
Adb11010110000	(	adb11010110000,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m010110_0	),
Adb11010110001	(	adb11010110001,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m010110_0	),
Adb11010110010	(	adb11010110010,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m010110_0	),
Adb11010110011	(	adb11010110011,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m010110_0	),
Adb11010110100	(	adb11010110100,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m010110_0	),
Adb11010110101	(	adb11010110101,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m010110_0	),
Adb11010110110	(	adb11010110110,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m010110_0	),
Adb11010110111	(	adb11010110111,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m010110_0	),
Adb11010111000	(	adb11010111000,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m010110_0	),
Adb11010111001	(	adb11010111001,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m010110_0	),
Adb11010111010	(	adb11010111010,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m010110_0	),
Adb11010111011	(	adb11010111011,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m010110_0	),
Adb11010111100	(	adb11010111100,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m010110_0	),
Adb11010111101	(	adb11010111101,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m010110_0	),
Adb11010111110	(	adb11010111110,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m010110_0	),
Adb11010111111	(	adb11010111111,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m010110_0	),
Adb11011000000	(	adb11011000000,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m010110_0	),
Adb11011000001	(	adb11011000001,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m010110_0	),
Adb11011000010	(	adb11011000010,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m010110_0	),
Adb11011000011	(	adb11011000011,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m010110_0	),
Adb11011000100	(	adb11011000100,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m010110_0	),
Adb11011000101	(	adb11011000101,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m010110_0	),
Adb11011000110	(	adb11011000110,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m010110_0	),
Adb11011000111	(	adb11011000111,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m010110_0	),
Adb11011001000	(	adb11011001000,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m010110_0	),
Adb11011001001	(	adb11011001001,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m010110_0	),
Adb11011001010	(	adb11011001010,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m010110_0	),
Adb11011001011	(	adb11011001011,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m010110_0	),
Adb11011001100	(	adb11011001100,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m010110_0	),
Adb11011001101	(	adb11011001101,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m010110_0	),
Adb11011001110	(	adb11011001110,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m010110_0	),
Adb11011001111	(	adb11011001111,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m010110_0	),
Adb11011010000	(	adb11011010000,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m010110_0	),
Adb11011010001	(	adb11011010001,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m010110_0	),
Adb11011010010	(	adb11011010010,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m010110_0	),
Adb11011010011	(	adb11011010011,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m010110_0	),
Adb11011010100	(	adb11011010100,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m010110_0	),
Adb11011010101	(	adb11011010101,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m010110_0	),
Adb11011010110	(	adb11011010110,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m010110_0	),
Adb11011010111	(	adb11011010111,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m010110_0	),
Adb11011011000	(	adb11011011000,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m010110_0	),
Adb11011011001	(	adb11011011001,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m010110_0	),
Adb11011011010	(	adb11011011010,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m010110_0	),
Adb11011011011	(	adb11011011011,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m010110_0	),
Adb11011011100	(	adb11011011100,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m010110_0	),
Adb11011011101	(	adb11011011101,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m010110_0	),
Adb11011011110	(	adb11011011110,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m010110_0	),
Adb11011011111	(	adb11011011111,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m010110_0	),
Adb11011100000	(	adb11011100000,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m010110_0	),
Adb11011100001	(	adb11011100001,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m010110_0	),
Adb11011100010	(	adb11011100010,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m010110_0	),
Adb11011100011	(	adb11011100011,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m010110_0	),
Adb11011100100	(	adb11011100100,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m010110_0	),
Adb11011100101	(	adb11011100101,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m010110_0	),
Adb11011100110	(	adb11011100110,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m010110_0	),
Adb11011100111	(	adb11011100111,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m010110_0	),
Adb11011101000	(	adb11011101000,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m010110_0	),
Adb11011101001	(	adb11011101001,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m010110_0	),
Adb11011101010	(	adb11011101010,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m010110_0	),
Adb11011101011	(	adb11011101011,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m010110_0	),
Adb11011101100	(	adb11011101100,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m010110_0	),
Adb11011101101	(	adb11011101101,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m010110_0	),
Adb11011101110	(	adb11011101110,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m010110_0	),
Adb11011101111	(	adb11011101111,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m010110_0	),
Adb11011110000	(	adb11011110000,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m010110_0	),
Adb11011110001	(	adb11011110001,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m010110_0	),
Adb11011110010	(	adb11011110010,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m010110_0	),
Adb11011110011	(	adb11011110011,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m010110_0	),
Adb11011110100	(	adb11011110100,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m010110_0	),
Adb11011110101	(	adb11011110101,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m010110_0	),
Adb11011110110	(	adb11011110110,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m010110_0	),
Adb11011110111	(	adb11011110111,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m010110_0	),
Adb11011111000	(	adb11011111000,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m010110_0	),
Adb11011111001	(	adb11011111001,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m010110_0	),
Adb11011111010	(	adb11011111010,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m010110_0	),
Adb11011111011	(	adb11011111011,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m010110_0	),
Adb11011111100	(	adb11011111100,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m010110_0	),
Adb11011111101	(	adb11011111101,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m010110_0	),
Adb11011111110	(	adb11011111110,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m010110_0	),
Adb11011111111	(	adb11011111111,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m010110_0	),
Adb11100000000	(	adb11100000000,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m001110_0	),
Adb11100000001	(	adb11100000001,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m001110_0	),
Adb11100000010	(	adb11100000010,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m001110_0	),
Adb11100000011	(	adb11100000011,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m001110_0	),
Adb11100000100	(	adb11100000100,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m001110_0	),
Adb11100000101	(	adb11100000101,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m001110_0	),
Adb11100000110	(	adb11100000110,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m001110_0	),
Adb11100000111	(	adb11100000111,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m001110_0	),
Adb11100001000	(	adb11100001000,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m001110_0	),
Adb11100001001	(	adb11100001001,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m001110_0	),
Adb11100001010	(	adb11100001010,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m001110_0	),
Adb11100001011	(	adb11100001011,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m001110_0	),
Adb11100001100	(	adb11100001100,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m001110_0	),
Adb11100001101	(	adb11100001101,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m001110_0	),
Adb11100001110	(	adb11100001110,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m001110_0	),
Adb11100001111	(	adb11100001111,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m001110_0	),
Adb11100010000	(	adb11100010000,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m001110_0	),
Adb11100010001	(	adb11100010001,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m001110_0	),
Adb11100010010	(	adb11100010010,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m001110_0	),
Adb11100010011	(	adb11100010011,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m001110_0	),
Adb11100010100	(	adb11100010100,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m001110_0	),
Adb11100010101	(	adb11100010101,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m001110_0	),
Adb11100010110	(	adb11100010110,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m001110_0	),
Adb11100010111	(	adb11100010111,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m001110_0	),
Adb11100011000	(	adb11100011000,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m001110_0	),
Adb11100011001	(	adb11100011001,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m001110_0	),
Adb11100011010	(	adb11100011010,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m001110_0	),
Adb11100011011	(	adb11100011011,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m001110_0	),
Adb11100011100	(	adb11100011100,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m001110_0	),
Adb11100011101	(	adb11100011101,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m001110_0	),
Adb11100011110	(	adb11100011110,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m001110_0	),
Adb11100011111	(	adb11100011111,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m001110_0	),
Adb11100100000	(	adb11100100000,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m001110_0	),
Adb11100100001	(	adb11100100001,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m001110_0	),
Adb11100100010	(	adb11100100010,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m001110_0	),
Adb11100100011	(	adb11100100011,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m001110_0	),
Adb11100100100	(	adb11100100100,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m001110_0	),
Adb11100100101	(	adb11100100101,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m001110_0	),
Adb11100100110	(	adb11100100110,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m001110_0	),
Adb11100100111	(	adb11100100111,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m001110_0	),
Adb11100101000	(	adb11100101000,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m001110_0	),
Adb11100101001	(	adb11100101001,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m001110_0	),
Adb11100101010	(	adb11100101010,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m001110_0	),
Adb11100101011	(	adb11100101011,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m001110_0	),
Adb11100101100	(	adb11100101100,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m001110_0	),
Adb11100101101	(	adb11100101101,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m001110_0	),
Adb11100101110	(	adb11100101110,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m001110_0	),
Adb11100101111	(	adb11100101111,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m001110_0	),
Adb11100110000	(	adb11100110000,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m001110_0	),
Adb11100110001	(	adb11100110001,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m001110_0	),
Adb11100110010	(	adb11100110010,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m001110_0	),
Adb11100110011	(	adb11100110011,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m001110_0	),
Adb11100110100	(	adb11100110100,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m001110_0	),
Adb11100110101	(	adb11100110101,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m001110_0	),
Adb11100110110	(	adb11100110110,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m001110_0	),
Adb11100110111	(	adb11100110111,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m001110_0	),
Adb11100111000	(	adb11100111000,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m001110_0	),
Adb11100111001	(	adb11100111001,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m001110_0	),
Adb11100111010	(	adb11100111010,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m001110_0	),
Adb11100111011	(	adb11100111011,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m001110_0	),
Adb11100111100	(	adb11100111100,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m001110_0	),
Adb11100111101	(	adb11100111101,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m001110_0	),
Adb11100111110	(	adb11100111110,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m001110_0	),
Adb11100111111	(	adb11100111111,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m001110_0	),
Adb11101000000	(	adb11101000000,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m001110_0	),
Adb11101000001	(	adb11101000001,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m001110_0	),
Adb11101000010	(	adb11101000010,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m001110_0	),
Adb11101000011	(	adb11101000011,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m001110_0	),
Adb11101000100	(	adb11101000100,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m001110_0	),
Adb11101000101	(	adb11101000101,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m001110_0	),
Adb11101000110	(	adb11101000110,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m001110_0	),
Adb11101000111	(	adb11101000111,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m001110_0	),
Adb11101001000	(	adb11101001000,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m001110_0	),
Adb11101001001	(	adb11101001001,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m001110_0	),
Adb11101001010	(	adb11101001010,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m001110_0	),
Adb11101001011	(	adb11101001011,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m001110_0	),
Adb11101001100	(	adb11101001100,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m001110_0	),
Adb11101001101	(	adb11101001101,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m001110_0	),
Adb11101001110	(	adb11101001110,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m001110_0	),
Adb11101001111	(	adb11101001111,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m001110_0	),
Adb11101010000	(	adb11101010000,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m001110_0	),
Adb11101010001	(	adb11101010001,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m001110_0	),
Adb11101010010	(	adb11101010010,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m001110_0	),
Adb11101010011	(	adb11101010011,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m001110_0	),
Adb11101010100	(	adb11101010100,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m001110_0	),
Adb11101010101	(	adb11101010101,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m001110_0	),
Adb11101010110	(	adb11101010110,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m001110_0	),
Adb11101010111	(	adb11101010111,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m001110_0	),
Adb11101011000	(	adb11101011000,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m001110_0	),
Adb11101011001	(	adb11101011001,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m001110_0	),
Adb11101011010	(	adb11101011010,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m001110_0	),
Adb11101011011	(	adb11101011011,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m001110_0	),
Adb11101011100	(	adb11101011100,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m001110_0	),
Adb11101011101	(	adb11101011101,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m001110_0	),
Adb11101011110	(	adb11101011110,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m001110_0	),
Adb11101011111	(	adb11101011111,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m001110_0	),
Adb11101100000	(	adb11101100000,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m001110_0	),
Adb11101100001	(	adb11101100001,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m001110_0	),
Adb11101100010	(	adb11101100010,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m001110_0	),
Adb11101100011	(	adb11101100011,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m001110_0	),
Adb11101100100	(	adb11101100100,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m001110_0	),
Adb11101100101	(	adb11101100101,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m001110_0	),
Adb11101100110	(	adb11101100110,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m001110_0	),
Adb11101100111	(	adb11101100111,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m001110_0	),
Adb11101101000	(	adb11101101000,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m001110_0	),
Adb11101101001	(	adb11101101001,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m001110_0	),
Adb11101101010	(	adb11101101010,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m001110_0	),
Adb11101101011	(	adb11101101011,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m001110_0	),
Adb11101101100	(	adb11101101100,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m001110_0	),
Adb11101101101	(	adb11101101101,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m001110_0	),
Adb11101101110	(	adb11101101110,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m001110_0	),
Adb11101101111	(	adb11101101111,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m001110_0	),
Adb11101110000	(	adb11101110000,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m001110_0	),
Adb11101110001	(	adb11101110001,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m001110_0	),
Adb11101110010	(	adb11101110010,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m001110_0	),
Adb11101110011	(	adb11101110011,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m001110_0	),
Adb11101110100	(	adb11101110100,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m001110_0	),
Adb11101110101	(	adb11101110101,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m001110_0	),
Adb11101110110	(	adb11101110110,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m001110_0	),
Adb11101110111	(	adb11101110111,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m001110_0	),
Adb11101111000	(	adb11101111000,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m001110_0	),
Adb11101111001	(	adb11101111001,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m001110_0	),
Adb11101111010	(	adb11101111010,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m001110_0	),
Adb11101111011	(	adb11101111011,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m001110_0	),
Adb11101111100	(	adb11101111100,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m001110_0	),
Adb11101111101	(	adb11101111101,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m001110_0	),
Adb11101111110	(	adb11101111110,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m001110_0	),
Adb11101111111	(	adb11101111111,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m001110_0	),
Adb11110000000	(	adb11110000000,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m000110_0	),
Adb11110000001	(	adb11110000001,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m000110_0	),
Adb11110000010	(	adb11110000010,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m000110_0	),
Adb11110000011	(	adb11110000011,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m000110_0	),
Adb11110000100	(	adb11110000100,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m000110_0	),
Adb11110000101	(	adb11110000101,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m000110_0	),
Adb11110000110	(	adb11110000110,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m000110_0	),
Adb11110000111	(	adb11110000111,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m000110_0	),
Adb11110001000	(	adb11110001000,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m000110_0	),
Adb11110001001	(	adb11110001001,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m000110_0	),
Adb11110001010	(	adb11110001010,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m000110_0	),
Adb11110001011	(	adb11110001011,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m000110_0	),
Adb11110001100	(	adb11110001100,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m000110_0	),
Adb11110001101	(	adb11110001101,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m000110_0	),
Adb11110001110	(	adb11110001110,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m000110_0	),
Adb11110001111	(	adb11110001111,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m000110_0	),
Adb11110010000	(	adb11110010000,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m000110_0	),
Adb11110010001	(	adb11110010001,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m000110_0	),
Adb11110010010	(	adb11110010010,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m000110_0	),
Adb11110010011	(	adb11110010011,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m000110_0	),
Adb11110010100	(	adb11110010100,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m000110_0	),
Adb11110010101	(	adb11110010101,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m000110_0	),
Adb11110010110	(	adb11110010110,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m000110_0	),
Adb11110010111	(	adb11110010111,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m000110_0	),
Adb11110011000	(	adb11110011000,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m000110_0	),
Adb11110011001	(	adb11110011001,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m000110_0	),
Adb11110011010	(	adb11110011010,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m000110_0	),
Adb11110011011	(	adb11110011011,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m000110_0	),
Adb11110011100	(	adb11110011100,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m000110_0	),
Adb11110011101	(	adb11110011101,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m000110_0	),
Adb11110011110	(	adb11110011110,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m000110_0	),
Adb11110011111	(	adb11110011111,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m000110_0	),
Adb11110100000	(	adb11110100000,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m000110_0	),
Adb11110100001	(	adb11110100001,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m000110_0	),
Adb11110100010	(	adb11110100010,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m000110_0	),
Adb11110100011	(	adb11110100011,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m000110_0	),
Adb11110100100	(	adb11110100100,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m000110_0	),
Adb11110100101	(	adb11110100101,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m000110_0	),
Adb11110100110	(	adb11110100110,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m000110_0	),
Adb11110100111	(	adb11110100111,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m000110_0	),
Adb11110101000	(	adb11110101000,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m000110_0	),
Adb11110101001	(	adb11110101001,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m000110_0	),
Adb11110101010	(	adb11110101010,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m000110_0	),
Adb11110101011	(	adb11110101011,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m000110_0	),
Adb11110101100	(	adb11110101100,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m000110_0	),
Adb11110101101	(	adb11110101101,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m000110_0	),
Adb11110101110	(	adb11110101110,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m000110_0	),
Adb11110101111	(	adb11110101111,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m000110_0	),
Adb11110110000	(	adb11110110000,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m000110_0	),
Adb11110110001	(	adb11110110001,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m000110_0	),
Adb11110110010	(	adb11110110010,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m000110_0	),
Adb11110110011	(	adb11110110011,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m000110_0	),
Adb11110110100	(	adb11110110100,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m000110_0	),
Adb11110110101	(	adb11110110101,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m000110_0	),
Adb11110110110	(	adb11110110110,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m000110_0	),
Adb11110110111	(	adb11110110111,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m000110_0	),
Adb11110111000	(	adb11110111000,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m000110_0	),
Adb11110111001	(	adb11110111001,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m000110_0	),
Adb11110111010	(	adb11110111010,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m000110_0	),
Adb11110111011	(	adb11110111011,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m000110_0	),
Adb11110111100	(	adb11110111100,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m000110_0	),
Adb11110111101	(	adb11110111101,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m000110_0	),
Adb11110111110	(	adb11110111110,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m000110_0	),
Adb11110111111	(	adb11110111111,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m000110_0	),
Adb11111000000	(	adb11111000000,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m000110_0	),
Adb11111000001	(	adb11111000001,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m000110_0	),
Adb11111000010	(	adb11111000010,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m000110_0	),
Adb11111000011	(	adb11111000011,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m000110_0	),
Adb11111000100	(	adb11111000100,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m000110_0	),
Adb11111000101	(	adb11111000101,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m000110_0	),
Adb11111000110	(	adb11111000110,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m000110_0	),
Adb11111000111	(	adb11111000111,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m000110_0	),
Adb11111001000	(	adb11111001000,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m000110_0	),
Adb11111001001	(	adb11111001001,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m000110_0	),
Adb11111001010	(	adb11111001010,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m000110_0	),
Adb11111001011	(	adb11111001011,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m000110_0	),
Adb11111001100	(	adb11111001100,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m000110_0	),
Adb11111001101	(	adb11111001101,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m000110_0	),
Adb11111001110	(	adb11111001110,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m000110_0	),
Adb11111001111	(	adb11111001111,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m000110_0	),
Adb11111010000	(	adb11111010000,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m000110_0	),
Adb11111010001	(	adb11111010001,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m000110_0	),
Adb11111010010	(	adb11111010010,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m000110_0	),
Adb11111010011	(	adb11111010011,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m000110_0	),
Adb11111010100	(	adb11111010100,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m000110_0	),
Adb11111010101	(	adb11111010101,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m000110_0	),
Adb11111010110	(	adb11111010110,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m000110_0	),
Adb11111010111	(	adb11111010111,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m000110_0	),
Adb11111011000	(	adb11111011000,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m000110_0	),
Adb11111011001	(	adb11111011001,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m000110_0	),
Adb11111011010	(	adb11111011010,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m000110_0	),
Adb11111011011	(	adb11111011011,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m000110_0	),
Adb11111011100	(	adb11111011100,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m000110_0	),
Adb11111011101	(	adb11111011101,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m000110_0	),
Adb11111011110	(	adb11111011110,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m000110_0	),
Adb11111011111	(	adb11111011111,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m000110_0	),
Adb11111100000	(	adb11111100000,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m000110_0	),
Adb11111100001	(	adb11111100001,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m000110_0	),
Adb11111100010	(	adb11111100010,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m000110_0	),
Adb11111100011	(	adb11111100011,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m000110_0	),
Adb11111100100	(	adb11111100100,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m000110_0	),
Adb11111100101	(	adb11111100101,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m000110_0	),
Adb11111100110	(	adb11111100110,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m000110_0	),
Adb11111100111	(	adb11111100111,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m000110_0	),
Adb11111101000	(	adb11111101000,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m000110_0	),
Adb11111101001	(	adb11111101001,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m000110_0	),
Adb11111101010	(	adb11111101010,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m000110_0	),
Adb11111101011	(	adb11111101011,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m000110_0	),
Adb11111101100	(	adb11111101100,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m000110_0	),
Adb11111101101	(	adb11111101101,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m000110_0	),
Adb11111101110	(	adb11111101110,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m000110_0	),
Adb11111101111	(	adb11111101111,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m000110_0	),
Adb11111110000	(	adb11111110000,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m000110_0	),
Adb11111110001	(	adb11111110001,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m000110_0	),
Adb11111110010	(	adb11111110010,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m000110_0	),
Adb11111110011	(	adb11111110011,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m000110_0	),
Adb11111110100	(	adb11111110100,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m000110_0	),
Adb11111110101	(	adb11111110101,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m000110_0	),
Adb11111110110	(	adb11111110110,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m000110_0	),
Adb11111110111	(	adb11111110111,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m000110_0	),
Adb11111111000	(	adb11111111000,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m000110_0	),
Adb11111111001	(	adb11111111001,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m000110_0	),
Adb11111111010	(	adb11111111010,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m000110_0	),
Adb11111111011	(	adb11111111011,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m000110_0	),
Adb11111111100	(	adb11111111100,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m000110_0	),
Adb11111111101	(	adb11111111101,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m000110_0	),
Adb11111111110	(	adb11111111110,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m000110_0	),
Adb11111111111	(	adb11111111111,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m000110_0	),
       Adb200(adb200,n0011,n0010,n0009,dbv1),
       Adb201(adb201,n0011,n0010,m0009,m0012),
       Adb210(adb210,n0011,m0010,n0009,m0019),
       Adb211(adb211,n0011,m0010,m0009,dbv0),
Adb20000000000	(	adb20000000000,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m111101_0	),
Adb20000000001	(	adb20000000001,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m111101_0	),
Adb20000000010	(	adb20000000010,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m111101_0	),
Adb20000000011	(	adb20000000011,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m111101_0	),
Adb20000000100	(	adb20000000100,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m111101_0	),
Adb20000000101	(	adb20000000101,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m111101_0	),
Adb20000000110	(	adb20000000110,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m111101_0	),
Adb20000000111	(	adb20000000111,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m111101_0	),
Adb20000001000	(	adb20000001000,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m111101_0	),
Adb20000001001	(	adb20000001001,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m111101_0	),
Adb20000001010	(	adb20000001010,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m111101_0	),
Adb20000001011	(	adb20000001011,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m111101_0	),
Adb20000001100	(	adb20000001100,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m111101_0	),
Adb20000001101	(	adb20000001101,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m111101_0	),
Adb20000001110	(	adb20000001110,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m111101_0	),
Adb20000001111	(	adb20000001111,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m111101_0	),
Adb20000010000	(	adb20000010000,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m111101_0	),
Adb20000010001	(	adb20000010001,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m111101_0	),
Adb20000010010	(	adb20000010010,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m111101_0	),
Adb20000010011	(	adb20000010011,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m111101_0	),
Adb20000010100	(	adb20000010100,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m111101_0	),
Adb20000010101	(	adb20000010101,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m111101_0	),
Adb20000010110	(	adb20000010110,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m111101_0	),
Adb20000010111	(	adb20000010111,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m111101_0	),
Adb20000011000	(	adb20000011000,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m111101_0	),
Adb20000011001	(	adb20000011001,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m111101_0	),
Adb20000011010	(	adb20000011010,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m111101_0	),
Adb20000011011	(	adb20000011011,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m111101_0	),
Adb20000011100	(	adb20000011100,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m111101_0	),
Adb20000011101	(	adb20000011101,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m111101_0	),
Adb20000011110	(	adb20000011110,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m111101_0	),
Adb20000011111	(	adb20000011111,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m111101_0	),
Adb20000100000	(	adb20000100000,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m111101_0	),
Adb20000100001	(	adb20000100001,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m111101_0	),
Adb20000100010	(	adb20000100010,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m111101_0	),
Adb20000100011	(	adb20000100011,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m111101_0	),
Adb20000100100	(	adb20000100100,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m111101_0	),
Adb20000100101	(	adb20000100101,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m111101_0	),
Adb20000100110	(	adb20000100110,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m111101_0	),
Adb20000100111	(	adb20000100111,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m111101_0	),
Adb20000101000	(	adb20000101000,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m111101_0	),
Adb20000101001	(	adb20000101001,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m111101_0	),
Adb20000101010	(	adb20000101010,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m111101_0	),
Adb20000101011	(	adb20000101011,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m111101_0	),
Adb20000101100	(	adb20000101100,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m111101_0	),
Adb20000101101	(	adb20000101101,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m111101_0	),
Adb20000101110	(	adb20000101110,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m111101_0	),
Adb20000101111	(	adb20000101111,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m111101_0	),
Adb20000110000	(	adb20000110000,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m111101_0	),
Adb20000110001	(	adb20000110001,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m111101_0	),
Adb20000110010	(	adb20000110010,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m111101_0	),
Adb20000110011	(	adb20000110011,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m111101_0	),
Adb20000110100	(	adb20000110100,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m111101_0	),
Adb20000110101	(	adb20000110101,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m111101_0	),
Adb20000110110	(	adb20000110110,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m111101_0	),
Adb20000110111	(	adb20000110111,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m111101_0	),
Adb20000111000	(	adb20000111000,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m111101_0	),
Adb20000111001	(	adb20000111001,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m111101_0	),
Adb20000111010	(	adb20000111010,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m111101_0	),
Adb20000111011	(	adb20000111011,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m111101_0	),
Adb20000111100	(	adb20000111100,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m111101_0	),
Adb20000111101	(	adb20000111101,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m111101_0	),
Adb20000111110	(	adb20000111110,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m111101_0	),
Adb20000111111	(	adb20000111111,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m111101_0	),
Adb20001000000	(	adb20001000000,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m111101_0	),
Adb20001000001	(	adb20001000001,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m111101_0	),
Adb20001000010	(	adb20001000010,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m111101_0	),
Adb20001000011	(	adb20001000011,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m111101_0	),
Adb20001000100	(	adb20001000100,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m111101_0	),
Adb20001000101	(	adb20001000101,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m111101_0	),
Adb20001000110	(	adb20001000110,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m111101_0	),
Adb20001000111	(	adb20001000111,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m111101_0	),
Adb20001001000	(	adb20001001000,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m111101_0	),
Adb20001001001	(	adb20001001001,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m111101_0	),
Adb20001001010	(	adb20001001010,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m111101_0	),
Adb20001001011	(	adb20001001011,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m111101_0	),
Adb20001001100	(	adb20001001100,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m111101_0	),
Adb20001001101	(	adb20001001101,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m111101_0	),
Adb20001001110	(	adb20001001110,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m111101_0	),
Adb20001001111	(	adb20001001111,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m111101_0	),
Adb20001010000	(	adb20001010000,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m111101_0	),
Adb20001010001	(	adb20001010001,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m111101_0	),
Adb20001010010	(	adb20001010010,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m111101_0	),
Adb20001010011	(	adb20001010011,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m111101_0	),
Adb20001010100	(	adb20001010100,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m111101_0	),
Adb20001010101	(	adb20001010101,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m111101_0	),
Adb20001010110	(	adb20001010110,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m111101_0	),
Adb20001010111	(	adb20001010111,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m111101_0	),
Adb20001011000	(	adb20001011000,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m111101_0	),
Adb20001011001	(	adb20001011001,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m111101_0	),
Adb20001011010	(	adb20001011010,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m111101_0	),
Adb20001011011	(	adb20001011011,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m111101_0	),
Adb20001011100	(	adb20001011100,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m111101_0	),
Adb20001011101	(	adb20001011101,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m111101_0	),
Adb20001011110	(	adb20001011110,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m111101_0	),
Adb20001011111	(	adb20001011111,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m111101_0	),
Adb20001100000	(	adb20001100000,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m111101_0	),
Adb20001100001	(	adb20001100001,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m111101_0	),
Adb20001100010	(	adb20001100010,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m111101_0	),
Adb20001100011	(	adb20001100011,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m111101_0	),
Adb20001100100	(	adb20001100100,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m111101_0	),
Adb20001100101	(	adb20001100101,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m111101_0	),
Adb20001100110	(	adb20001100110,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m111101_0	),
Adb20001100111	(	adb20001100111,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m111101_0	),
Adb20001101000	(	adb20001101000,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m111101_0	),
Adb20001101001	(	adb20001101001,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m111101_0	),
Adb20001101010	(	adb20001101010,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m111101_0	),
Adb20001101011	(	adb20001101011,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m111101_0	),
Adb20001101100	(	adb20001101100,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m111101_0	),
Adb20001101101	(	adb20001101101,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m111101_0	),
Adb20001101110	(	adb20001101110,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m111101_0	),
Adb20001101111	(	adb20001101111,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m111101_0	),
Adb20001110000	(	adb20001110000,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m111101_0	),
Adb20001110001	(	adb20001110001,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m111101_0	),
Adb20001110010	(	adb20001110010,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m111101_0	),
Adb20001110011	(	adb20001110011,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m111101_0	),
Adb20001110100	(	adb20001110100,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m111101_0	),
Adb20001110101	(	adb20001110101,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m111101_0	),
Adb20001110110	(	adb20001110110,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m111101_0	),
Adb20001110111	(	adb20001110111,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m111101_0	),
Adb20001111000	(	adb20001111000,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m111101_0	),
Adb20001111001	(	adb20001111001,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m111101_0	),
Adb20001111010	(	adb20001111010,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m111101_0	),
Adb20001111011	(	adb20001111011,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m111101_0	),
Adb20001111100	(	adb20001111100,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m111101_0	),
Adb20001111101	(	adb20001111101,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m111101_0	),
Adb20001111110	(	adb20001111110,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m111101_0	),
Adb20001111111	(	adb20001111111,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m111101_0	),
Adb20010000000	(	adb20010000000,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m110101_0	),
Adb20010000001	(	adb20010000001,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m110101_0	),
Adb20010000010	(	adb20010000010,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m110101_0	),
Adb20010000011	(	adb20010000011,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m110101_0	),
Adb20010000100	(	adb20010000100,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m110101_0	),
Adb20010000101	(	adb20010000101,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m110101_0	),
Adb20010000110	(	adb20010000110,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m110101_0	),
Adb20010000111	(	adb20010000111,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m110101_0	),
Adb20010001000	(	adb20010001000,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m110101_0	),
Adb20010001001	(	adb20010001001,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m110101_0	),
Adb20010001010	(	adb20010001010,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m110101_0	),
Adb20010001011	(	adb20010001011,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m110101_0	),
Adb20010001100	(	adb20010001100,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m110101_0	),
Adb20010001101	(	adb20010001101,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m110101_0	),
Adb20010001110	(	adb20010001110,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m110101_0	),
Adb20010001111	(	adb20010001111,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m110101_0	),
Adb20010010000	(	adb20010010000,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m110101_0	),
Adb20010010001	(	adb20010010001,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m110101_0	),
Adb20010010010	(	adb20010010010,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m110101_0	),
Adb20010010011	(	adb20010010011,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m110101_0	),
Adb20010010100	(	adb20010010100,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m110101_0	),
Adb20010010101	(	adb20010010101,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m110101_0	),
Adb20010010110	(	adb20010010110,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m110101_0	),
Adb20010010111	(	adb20010010111,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m110101_0	),
Adb20010011000	(	adb20010011000,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m110101_0	),
Adb20010011001	(	adb20010011001,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m110101_0	),
Adb20010011010	(	adb20010011010,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m110101_0	),
Adb20010011011	(	adb20010011011,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m110101_0	),
Adb20010011100	(	adb20010011100,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m110101_0	),
Adb20010011101	(	adb20010011101,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m110101_0	),
Adb20010011110	(	adb20010011110,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m110101_0	),
Adb20010011111	(	adb20010011111,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m110101_0	),
Adb20010100000	(	adb20010100000,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m110101_0	),
Adb20010100001	(	adb20010100001,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m110101_0	),
Adb20010100010	(	adb20010100010,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m110101_0	),
Adb20010100011	(	adb20010100011,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m110101_0	),
Adb20010100100	(	adb20010100100,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m110101_0	),
Adb20010100101	(	adb20010100101,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m110101_0	),
Adb20010100110	(	adb20010100110,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m110101_0	),
Adb20010100111	(	adb20010100111,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m110101_0	),
Adb20010101000	(	adb20010101000,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m110101_0	),
Adb20010101001	(	adb20010101001,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m110101_0	),
Adb20010101010	(	adb20010101010,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m110101_0	),
Adb20010101011	(	adb20010101011,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m110101_0	),
Adb20010101100	(	adb20010101100,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m110101_0	),
Adb20010101101	(	adb20010101101,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m110101_0	),
Adb20010101110	(	adb20010101110,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m110101_0	),
Adb20010101111	(	adb20010101111,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m110101_0	),
Adb20010110000	(	adb20010110000,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m110101_0	),
Adb20010110001	(	adb20010110001,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m110101_0	),
Adb20010110010	(	adb20010110010,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m110101_0	),
Adb20010110011	(	adb20010110011,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m110101_0	),
Adb20010110100	(	adb20010110100,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m110101_0	),
Adb20010110101	(	adb20010110101,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m110101_0	),
Adb20010110110	(	adb20010110110,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m110101_0	),
Adb20010110111	(	adb20010110111,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m110101_0	),
Adb20010111000	(	adb20010111000,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m110101_0	),
Adb20010111001	(	adb20010111001,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m110101_0	),
Adb20010111010	(	adb20010111010,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m110101_0	),
Adb20010111011	(	adb20010111011,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m110101_0	),
Adb20010111100	(	adb20010111100,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m110101_0	),
Adb20010111101	(	adb20010111101,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m110101_0	),
Adb20010111110	(	adb20010111110,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m110101_0	),
Adb20010111111	(	adb20010111111,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m110101_0	),
Adb20011000000	(	adb20011000000,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m110101_0	),
Adb20011000001	(	adb20011000001,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m110101_0	),
Adb20011000010	(	adb20011000010,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m110101_0	),
Adb20011000011	(	adb20011000011,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m110101_0	),
Adb20011000100	(	adb20011000100,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m110101_0	),
Adb20011000101	(	adb20011000101,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m110101_0	),
Adb20011000110	(	adb20011000110,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m110101_0	),
Adb20011000111	(	adb20011000111,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m110101_0	),
Adb20011001000	(	adb20011001000,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m110101_0	),
Adb20011001001	(	adb20011001001,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m110101_0	),
Adb20011001010	(	adb20011001010,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m110101_0	),
Adb20011001011	(	adb20011001011,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m110101_0	),
Adb20011001100	(	adb20011001100,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m110101_0	),
Adb20011001101	(	adb20011001101,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m110101_0	),
Adb20011001110	(	adb20011001110,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m110101_0	),
Adb20011001111	(	adb20011001111,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m110101_0	),
Adb20011010000	(	adb20011010000,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m110101_0	),
Adb20011010001	(	adb20011010001,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m110101_0	),
Adb20011010010	(	adb20011010010,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m110101_0	),
Adb20011010011	(	adb20011010011,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m110101_0	),
Adb20011010100	(	adb20011010100,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m110101_0	),
Adb20011010101	(	adb20011010101,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m110101_0	),
Adb20011010110	(	adb20011010110,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m110101_0	),
Adb20011010111	(	adb20011010111,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m110101_0	),
Adb20011011000	(	adb20011011000,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m110101_0	),
Adb20011011001	(	adb20011011001,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m110101_0	),
Adb20011011010	(	adb20011011010,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m110101_0	),
Adb20011011011	(	adb20011011011,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m110101_0	),
Adb20011011100	(	adb20011011100,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m110101_0	),
Adb20011011101	(	adb20011011101,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m110101_0	),
Adb20011011110	(	adb20011011110,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m110101_0	),
Adb20011011111	(	adb20011011111,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m110101_0	),
Adb20011100000	(	adb20011100000,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m110101_0	),
Adb20011100001	(	adb20011100001,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m110101_0	),
Adb20011100010	(	adb20011100010,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m110101_0	),
Adb20011100011	(	adb20011100011,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m110101_0	),
Adb20011100100	(	adb20011100100,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m110101_0	),
Adb20011100101	(	adb20011100101,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m110101_0	),
Adb20011100110	(	adb20011100110,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m110101_0	),
Adb20011100111	(	adb20011100111,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m110101_0	),
Adb20011101000	(	adb20011101000,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m110101_0	),
Adb20011101001	(	adb20011101001,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m110101_0	),
Adb20011101010	(	adb20011101010,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m110101_0	),
Adb20011101011	(	adb20011101011,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m110101_0	),
Adb20011101100	(	adb20011101100,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m110101_0	),
Adb20011101101	(	adb20011101101,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m110101_0	),
Adb20011101110	(	adb20011101110,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m110101_0	),
Adb20011101111	(	adb20011101111,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m110101_0	),
Adb20011110000	(	adb20011110000,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m110101_0	),
Adb20011110001	(	adb20011110001,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m110101_0	),
Adb20011110010	(	adb20011110010,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m110101_0	),
Adb20011110011	(	adb20011110011,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m110101_0	),
Adb20011110100	(	adb20011110100,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m110101_0	),
Adb20011110101	(	adb20011110101,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m110101_0	),
Adb20011110110	(	adb20011110110,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m110101_0	),
Adb20011110111	(	adb20011110111,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m110101_0	),
Adb20011111000	(	adb20011111000,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m110101_0	),
Adb20011111001	(	adb20011111001,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m110101_0	),
Adb20011111010	(	adb20011111010,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m110101_0	),
Adb20011111011	(	adb20011111011,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m110101_0	),
Adb20011111100	(	adb20011111100,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m110101_0	),
Adb20011111101	(	adb20011111101,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m110101_0	),
Adb20011111110	(	adb20011111110,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m110101_0	),
Adb20011111111	(	adb20011111111,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m110101_0	),
Adb20100000000	(	adb20100000000,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m101101_0	),
Adb20100000001	(	adb20100000001,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m101101_0	),
Adb20100000010	(	adb20100000010,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m101101_0	),
Adb20100000011	(	adb20100000011,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m101101_0	),
Adb20100000100	(	adb20100000100,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m101101_0	),
Adb20100000101	(	adb20100000101,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m101101_0	),
Adb20100000110	(	adb20100000110,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m101101_0	),
Adb20100000111	(	adb20100000111,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m101101_0	),
Adb20100001000	(	adb20100001000,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m101101_0	),
Adb20100001001	(	adb20100001001,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m101101_0	),
Adb20100001010	(	adb20100001010,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m101101_0	),
Adb20100001011	(	adb20100001011,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m101101_0	),
Adb20100001100	(	adb20100001100,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m101101_0	),
Adb20100001101	(	adb20100001101,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m101101_0	),
Adb20100001110	(	adb20100001110,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m101101_0	),
Adb20100001111	(	adb20100001111,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m101101_0	),
Adb20100010000	(	adb20100010000,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m101101_0	),
Adb20100010001	(	adb20100010001,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m101101_0	),
Adb20100010010	(	adb20100010010,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m101101_0	),
Adb20100010011	(	adb20100010011,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m101101_0	),
Adb20100010100	(	adb20100010100,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m101101_0	),
Adb20100010101	(	adb20100010101,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m101101_0	),
Adb20100010110	(	adb20100010110,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m101101_0	),
Adb20100010111	(	adb20100010111,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m101101_0	),
Adb20100011000	(	adb20100011000,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m101101_0	),
Adb20100011001	(	adb20100011001,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m101101_0	),
Adb20100011010	(	adb20100011010,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m101101_0	),
Adb20100011011	(	adb20100011011,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m101101_0	),
Adb20100011100	(	adb20100011100,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m101101_0	),
Adb20100011101	(	adb20100011101,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m101101_0	),
Adb20100011110	(	adb20100011110,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m101101_0	),
Adb20100011111	(	adb20100011111,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m101101_0	),
Adb20100100000	(	adb20100100000,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m101101_0	),
Adb20100100001	(	adb20100100001,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m101101_0	),
Adb20100100010	(	adb20100100010,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m101101_0	),
Adb20100100011	(	adb20100100011,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m101101_0	),
Adb20100100100	(	adb20100100100,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m101101_0	),
Adb20100100101	(	adb20100100101,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m101101_0	),
Adb20100100110	(	adb20100100110,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m101101_0	),
Adb20100100111	(	adb20100100111,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m101101_0	),
Adb20100101000	(	adb20100101000,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m101101_0	),
Adb20100101001	(	adb20100101001,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m101101_0	),
Adb20100101010	(	adb20100101010,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m101101_0	),
Adb20100101011	(	adb20100101011,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m101101_0	),
Adb20100101100	(	adb20100101100,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m101101_0	),
Adb20100101101	(	adb20100101101,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m101101_0	),
Adb20100101110	(	adb20100101110,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m101101_0	),
Adb20100101111	(	adb20100101111,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m101101_0	),
Adb20100110000	(	adb20100110000,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m101101_0	),
Adb20100110001	(	adb20100110001,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m101101_0	),
Adb20100110010	(	adb20100110010,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m101101_0	),
Adb20100110011	(	adb20100110011,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m101101_0	),
Adb20100110100	(	adb20100110100,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m101101_0	),
Adb20100110101	(	adb20100110101,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m101101_0	),
Adb20100110110	(	adb20100110110,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m101101_0	),
Adb20100110111	(	adb20100110111,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m101101_0	),
Adb20100111000	(	adb20100111000,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m101101_0	),
Adb20100111001	(	adb20100111001,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m101101_0	),
Adb20100111010	(	adb20100111010,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m101101_0	),
Adb20100111011	(	adb20100111011,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m101101_0	),
Adb20100111100	(	adb20100111100,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m101101_0	),
Adb20100111101	(	adb20100111101,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m101101_0	),
Adb20100111110	(	adb20100111110,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m101101_0	),
Adb20100111111	(	adb20100111111,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m101101_0	),
Adb20101000000	(	adb20101000000,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m101101_0	),
Adb20101000001	(	adb20101000001,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m101101_0	),
Adb20101000010	(	adb20101000010,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m101101_0	),
Adb20101000011	(	adb20101000011,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m101101_0	),
Adb20101000100	(	adb20101000100,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m101101_0	),
Adb20101000101	(	adb20101000101,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m101101_0	),
Adb20101000110	(	adb20101000110,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m101101_0	),
Adb20101000111	(	adb20101000111,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m101101_0	),
Adb20101001000	(	adb20101001000,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m101101_0	),
Adb20101001001	(	adb20101001001,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m101101_0	),
Adb20101001010	(	adb20101001010,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m101101_0	),
Adb20101001011	(	adb20101001011,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m101101_0	),
Adb20101001100	(	adb20101001100,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m101101_0	),
Adb20101001101	(	adb20101001101,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m101101_0	),
Adb20101001110	(	adb20101001110,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m101101_0	),
Adb20101001111	(	adb20101001111,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m101101_0	),
Adb20101010000	(	adb20101010000,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m101101_0	),
Adb20101010001	(	adb20101010001,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m101101_0	),
Adb20101010010	(	adb20101010010,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m101101_0	),
Adb20101010011	(	adb20101010011,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m101101_0	),
Adb20101010100	(	adb20101010100,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m101101_0	),
Adb20101010101	(	adb20101010101,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m101101_0	),
Adb20101010110	(	adb20101010110,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m101101_0	),
Adb20101010111	(	adb20101010111,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m101101_0	),
Adb20101011000	(	adb20101011000,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m101101_0	),
Adb20101011001	(	adb20101011001,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m101101_0	),
Adb20101011010	(	adb20101011010,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m101101_0	),
Adb20101011011	(	adb20101011011,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m101101_0	),
Adb20101011100	(	adb20101011100,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m101101_0	),
Adb20101011101	(	adb20101011101,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m101101_0	),
Adb20101011110	(	adb20101011110,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m101101_0	),
Adb20101011111	(	adb20101011111,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m101101_0	),
Adb20101100000	(	adb20101100000,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m101101_0	),
Adb20101100001	(	adb20101100001,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m101101_0	),
Adb20101100010	(	adb20101100010,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m101101_0	),
Adb20101100011	(	adb20101100011,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m101101_0	),
Adb20101100100	(	adb20101100100,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m101101_0	),
Adb20101100101	(	adb20101100101,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m101101_0	),
Adb20101100110	(	adb20101100110,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m101101_0	),
Adb20101100111	(	adb20101100111,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m101101_0	),
Adb20101101000	(	adb20101101000,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m101101_0	),
Adb20101101001	(	adb20101101001,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m101101_0	),
Adb20101101010	(	adb20101101010,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m101101_0	),
Adb20101101011	(	adb20101101011,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m101101_0	),
Adb20101101100	(	adb20101101100,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m101101_0	),
Adb20101101101	(	adb20101101101,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m101101_0	),
Adb20101101110	(	adb20101101110,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m101101_0	),
Adb20101101111	(	adb20101101111,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m101101_0	),
Adb20101110000	(	adb20101110000,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m101101_0	),
Adb20101110001	(	adb20101110001,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m101101_0	),
Adb20101110010	(	adb20101110010,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m101101_0	),
Adb20101110011	(	adb20101110011,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m101101_0	),
Adb20101110100	(	adb20101110100,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m101101_0	),
Adb20101110101	(	adb20101110101,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m101101_0	),
Adb20101110110	(	adb20101110110,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m101101_0	),
Adb20101110111	(	adb20101110111,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m101101_0	),
Adb20101111000	(	adb20101111000,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m101101_0	),
Adb20101111001	(	adb20101111001,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m101101_0	),
Adb20101111010	(	adb20101111010,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m101101_0	),
Adb20101111011	(	adb20101111011,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m101101_0	),
Adb20101111100	(	adb20101111100,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m101101_0	),
Adb20101111101	(	adb20101111101,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m101101_0	),
Adb20101111110	(	adb20101111110,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m101101_0	),
Adb20101111111	(	adb20101111111,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m101101_0	),
Adb20110000000	(	adb20110000000,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m100101_0	),
Adb20110000001	(	adb20110000001,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m100101_0	),
Adb20110000010	(	adb20110000010,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m100101_0	),
Adb20110000011	(	adb20110000011,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m100101_0	),
Adb20110000100	(	adb20110000100,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m100101_0	),
Adb20110000101	(	adb20110000101,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m100101_0	),
Adb20110000110	(	adb20110000110,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m100101_0	),
Adb20110000111	(	adb20110000111,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m100101_0	),
Adb20110001000	(	adb20110001000,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m100101_0	),
Adb20110001001	(	adb20110001001,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m100101_0	),
Adb20110001010	(	adb20110001010,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m100101_0	),
Adb20110001011	(	adb20110001011,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m100101_0	),
Adb20110001100	(	adb20110001100,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m100101_0	),
Adb20110001101	(	adb20110001101,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m100101_0	),
Adb20110001110	(	adb20110001110,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m100101_0	),
Adb20110001111	(	adb20110001111,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m100101_0	),
Adb20110010000	(	adb20110010000,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m100101_0	),
Adb20110010001	(	adb20110010001,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m100101_0	),
Adb20110010010	(	adb20110010010,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m100101_0	),
Adb20110010011	(	adb20110010011,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m100101_0	),
Adb20110010100	(	adb20110010100,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m100101_0	),
Adb20110010101	(	adb20110010101,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m100101_0	),
Adb20110010110	(	adb20110010110,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m100101_0	),
Adb20110010111	(	adb20110010111,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m100101_0	),
Adb20110011000	(	adb20110011000,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m100101_0	),
Adb20110011001	(	adb20110011001,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m100101_0	),
Adb20110011010	(	adb20110011010,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m100101_0	),
Adb20110011011	(	adb20110011011,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m100101_0	),
Adb20110011100	(	adb20110011100,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m100101_0	),
Adb20110011101	(	adb20110011101,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m100101_0	),
Adb20110011110	(	adb20110011110,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m100101_0	),
Adb20110011111	(	adb20110011111,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m100101_0	),
Adb20110100000	(	adb20110100000,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m100101_0	),
Adb20110100001	(	adb20110100001,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m100101_0	),
Adb20110100010	(	adb20110100010,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m100101_0	),
Adb20110100011	(	adb20110100011,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m100101_0	),
Adb20110100100	(	adb20110100100,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m100101_0	),
Adb20110100101	(	adb20110100101,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m100101_0	),
Adb20110100110	(	adb20110100110,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m100101_0	),
Adb20110100111	(	adb20110100111,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m100101_0	),
Adb20110101000	(	adb20110101000,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m100101_0	),
Adb20110101001	(	adb20110101001,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m100101_0	),
Adb20110101010	(	adb20110101010,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m100101_0	),
Adb20110101011	(	adb20110101011,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m100101_0	),
Adb20110101100	(	adb20110101100,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m100101_0	),
Adb20110101101	(	adb20110101101,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m100101_0	),
Adb20110101110	(	adb20110101110,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m100101_0	),
Adb20110101111	(	adb20110101111,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m100101_0	),
Adb20110110000	(	adb20110110000,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m100101_0	),
Adb20110110001	(	adb20110110001,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m100101_0	),
Adb20110110010	(	adb20110110010,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m100101_0	),
Adb20110110011	(	adb20110110011,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m100101_0	),
Adb20110110100	(	adb20110110100,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m100101_0	),
Adb20110110101	(	adb20110110101,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m100101_0	),
Adb20110110110	(	adb20110110110,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m100101_0	),
Adb20110110111	(	adb20110110111,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m100101_0	),
Adb20110111000	(	adb20110111000,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m100101_0	),
Adb20110111001	(	adb20110111001,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m100101_0	),
Adb20110111010	(	adb20110111010,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m100101_0	),
Adb20110111011	(	adb20110111011,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m100101_0	),
Adb20110111100	(	adb20110111100,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m100101_0	),
Adb20110111101	(	adb20110111101,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m100101_0	),
Adb20110111110	(	adb20110111110,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m100101_0	),
Adb20110111111	(	adb20110111111,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m100101_0	),
Adb20111000000	(	adb20111000000,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m100101_0	),
Adb20111000001	(	adb20111000001,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m100101_0	),
Adb20111000010	(	adb20111000010,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m100101_0	),
Adb20111000011	(	adb20111000011,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m100101_0	),
Adb20111000100	(	adb20111000100,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m100101_0	),
Adb20111000101	(	adb20111000101,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m100101_0	),
Adb20111000110	(	adb20111000110,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m100101_0	),
Adb20111000111	(	adb20111000111,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m100101_0	),
Adb20111001000	(	adb20111001000,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m100101_0	),
Adb20111001001	(	adb20111001001,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m100101_0	),
Adb20111001010	(	adb20111001010,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m100101_0	),
Adb20111001011	(	adb20111001011,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m100101_0	),
Adb20111001100	(	adb20111001100,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m100101_0	),
Adb20111001101	(	adb20111001101,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m100101_0	),
Adb20111001110	(	adb20111001110,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m100101_0	),
Adb20111001111	(	adb20111001111,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m100101_0	),
Adb20111010000	(	adb20111010000,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m100101_0	),
Adb20111010001	(	adb20111010001,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m100101_0	),
Adb20111010010	(	adb20111010010,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m100101_0	),
Adb20111010011	(	adb20111010011,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m100101_0	),
Adb20111010100	(	adb20111010100,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m100101_0	),
Adb20111010101	(	adb20111010101,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m100101_0	),
Adb20111010110	(	adb20111010110,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m100101_0	),
Adb20111010111	(	adb20111010111,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m100101_0	),
Adb20111011000	(	adb20111011000,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m100101_0	),
Adb20111011001	(	adb20111011001,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m100101_0	),
Adb20111011010	(	adb20111011010,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m100101_0	),
Adb20111011011	(	adb20111011011,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m100101_0	),
Adb20111011100	(	adb20111011100,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m100101_0	),
Adb20111011101	(	adb20111011101,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m100101_0	),
Adb20111011110	(	adb20111011110,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m100101_0	),
Adb20111011111	(	adb20111011111,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m100101_0	),
Adb20111100000	(	adb20111100000,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m100101_0	),
Adb20111100001	(	adb20111100001,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m100101_0	),
Adb20111100010	(	adb20111100010,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m100101_0	),
Adb20111100011	(	adb20111100011,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m100101_0	),
Adb20111100100	(	adb20111100100,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m100101_0	),
Adb20111100101	(	adb20111100101,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m100101_0	),
Adb20111100110	(	adb20111100110,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m100101_0	),
Adb20111100111	(	adb20111100111,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m100101_0	),
Adb20111101000	(	adb20111101000,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m100101_0	),
Adb20111101001	(	adb20111101001,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m100101_0	),
Adb20111101010	(	adb20111101010,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m100101_0	),
Adb20111101011	(	adb20111101011,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m100101_0	),
Adb20111101100	(	adb20111101100,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m100101_0	),
Adb20111101101	(	adb20111101101,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m100101_0	),
Adb20111101110	(	adb20111101110,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m100101_0	),
Adb20111101111	(	adb20111101111,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m100101_0	),
Adb20111110000	(	adb20111110000,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m100101_0	),
Adb20111110001	(	adb20111110001,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m100101_0	),
Adb20111110010	(	adb20111110010,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m100101_0	),
Adb20111110011	(	adb20111110011,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m100101_0	),
Adb20111110100	(	adb20111110100,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m100101_0	),
Adb20111110101	(	adb20111110101,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m100101_0	),
Adb20111110110	(	adb20111110110,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m100101_0	),
Adb20111110111	(	adb20111110111,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m100101_0	),
Adb20111111000	(	adb20111111000,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m100101_0	),
Adb20111111001	(	adb20111111001,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m100101_0	),
Adb20111111010	(	adb20111111010,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m100101_0	),
Adb20111111011	(	adb20111111011,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m100101_0	),
Adb20111111100	(	adb20111111100,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m100101_0	),
Adb20111111101	(	adb20111111101,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m100101_0	),
Adb20111111110	(	adb20111111110,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m100101_0	),
Adb20111111111	(	adb20111111111,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m100101_0	),
Adb21000000000	(	adb21000000000,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m011101_0	),
Adb21000000001	(	adb21000000001,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m011101_0	),
Adb21000000010	(	adb21000000010,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m011101_0	),
Adb21000000011	(	adb21000000011,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m011101_0	),
Adb21000000100	(	adb21000000100,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m011101_0	),
Adb21000000101	(	adb21000000101,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m011101_0	),
Adb21000000110	(	adb21000000110,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m011101_0	),
Adb21000000111	(	adb21000000111,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m011101_0	),
Adb21000001000	(	adb21000001000,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m011101_0	),
Adb21000001001	(	adb21000001001,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m011101_0	),
Adb21000001010	(	adb21000001010,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m011101_0	),
Adb21000001011	(	adb21000001011,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m011101_0	),
Adb21000001100	(	adb21000001100,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m011101_0	),
Adb21000001101	(	adb21000001101,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m011101_0	),
Adb21000001110	(	adb21000001110,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m011101_0	),
Adb21000001111	(	adb21000001111,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m011101_0	),
Adb21000010000	(	adb21000010000,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m011101_0	),
Adb21000010001	(	adb21000010001,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m011101_0	),
Adb21000010010	(	adb21000010010,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m011101_0	),
Adb21000010011	(	adb21000010011,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m011101_0	),
Adb21000010100	(	adb21000010100,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m011101_0	),
Adb21000010101	(	adb21000010101,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m011101_0	),
Adb21000010110	(	adb21000010110,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m011101_0	),
Adb21000010111	(	adb21000010111,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m011101_0	),
Adb21000011000	(	adb21000011000,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m011101_0	),
Adb21000011001	(	adb21000011001,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m011101_0	),
Adb21000011010	(	adb21000011010,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m011101_0	),
Adb21000011011	(	adb21000011011,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m011101_0	),
Adb21000011100	(	adb21000011100,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m011101_0	),
Adb21000011101	(	adb21000011101,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m011101_0	),
Adb21000011110	(	adb21000011110,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m011101_0	),
Adb21000011111	(	adb21000011111,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m011101_0	),
Adb21000100000	(	adb21000100000,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m011101_0	),
Adb21000100001	(	adb21000100001,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m011101_0	),
Adb21000100010	(	adb21000100010,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m011101_0	),
Adb21000100011	(	adb21000100011,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m011101_0	),
Adb21000100100	(	adb21000100100,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m011101_0	),
Adb21000100101	(	adb21000100101,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m011101_0	),
Adb21000100110	(	adb21000100110,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m011101_0	),
Adb21000100111	(	adb21000100111,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m011101_0	),
Adb21000101000	(	adb21000101000,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m011101_0	),
Adb21000101001	(	adb21000101001,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m011101_0	),
Adb21000101010	(	adb21000101010,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m011101_0	),
Adb21000101011	(	adb21000101011,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m011101_0	),
Adb21000101100	(	adb21000101100,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m011101_0	),
Adb21000101101	(	adb21000101101,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m011101_0	),
Adb21000101110	(	adb21000101110,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m011101_0	),
Adb21000101111	(	adb21000101111,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m011101_0	),
Adb21000110000	(	adb21000110000,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m011101_0	),
Adb21000110001	(	adb21000110001,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m011101_0	),
Adb21000110010	(	adb21000110010,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m011101_0	),
Adb21000110011	(	adb21000110011,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m011101_0	),
Adb21000110100	(	adb21000110100,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m011101_0	),
Adb21000110101	(	adb21000110101,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m011101_0	),
Adb21000110110	(	adb21000110110,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m011101_0	),
Adb21000110111	(	adb21000110111,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m011101_0	),
Adb21000111000	(	adb21000111000,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m011101_0	),
Adb21000111001	(	adb21000111001,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m011101_0	),
Adb21000111010	(	adb21000111010,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m011101_0	),
Adb21000111011	(	adb21000111011,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m011101_0	),
Adb21000111100	(	adb21000111100,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m011101_0	),
Adb21000111101	(	adb21000111101,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m011101_0	),
Adb21000111110	(	adb21000111110,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m011101_0	),
Adb21000111111	(	adb21000111111,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m011101_0	),
Adb21001000000	(	adb21001000000,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m011101_0	),
Adb21001000001	(	adb21001000001,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m011101_0	),
Adb21001000010	(	adb21001000010,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m011101_0	),
Adb21001000011	(	adb21001000011,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m011101_0	),
Adb21001000100	(	adb21001000100,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m011101_0	),
Adb21001000101	(	adb21001000101,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m011101_0	),
Adb21001000110	(	adb21001000110,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m011101_0	),
Adb21001000111	(	adb21001000111,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m011101_0	),
Adb21001001000	(	adb21001001000,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m011101_0	),
Adb21001001001	(	adb21001001001,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m011101_0	),
Adb21001001010	(	adb21001001010,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m011101_0	),
Adb21001001011	(	adb21001001011,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m011101_0	),
Adb21001001100	(	adb21001001100,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m011101_0	),
Adb21001001101	(	adb21001001101,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m011101_0	),
Adb21001001110	(	adb21001001110,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m011101_0	),
Adb21001001111	(	adb21001001111,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m011101_0	),
Adb21001010000	(	adb21001010000,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m011101_0	),
Adb21001010001	(	adb21001010001,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m011101_0	),
Adb21001010010	(	adb21001010010,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m011101_0	),
Adb21001010011	(	adb21001010011,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m011101_0	),
Adb21001010100	(	adb21001010100,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m011101_0	),
Adb21001010101	(	adb21001010101,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m011101_0	),
Adb21001010110	(	adb21001010110,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m011101_0	),
Adb21001010111	(	adb21001010111,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m011101_0	),
Adb21001011000	(	adb21001011000,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m011101_0	),
Adb21001011001	(	adb21001011001,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m011101_0	),
Adb21001011010	(	adb21001011010,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m011101_0	),
Adb21001011011	(	adb21001011011,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m011101_0	),
Adb21001011100	(	adb21001011100,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m011101_0	),
Adb21001011101	(	adb21001011101,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m011101_0	),
Adb21001011110	(	adb21001011110,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m011101_0	),
Adb21001011111	(	adb21001011111,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m011101_0	),
Adb21001100000	(	adb21001100000,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m011101_0	),
Adb21001100001	(	adb21001100001,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m011101_0	),
Adb21001100010	(	adb21001100010,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m011101_0	),
Adb21001100011	(	adb21001100011,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m011101_0	),
Adb21001100100	(	adb21001100100,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m011101_0	),
Adb21001100101	(	adb21001100101,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m011101_0	),
Adb21001100110	(	adb21001100110,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m011101_0	),
Adb21001100111	(	adb21001100111,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m011101_0	),
Adb21001101000	(	adb21001101000,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m011101_0	),
Adb21001101001	(	adb21001101001,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m011101_0	),
Adb21001101010	(	adb21001101010,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m011101_0	),
Adb21001101011	(	adb21001101011,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m011101_0	),
Adb21001101100	(	adb21001101100,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m011101_0	),
Adb21001101101	(	adb21001101101,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m011101_0	),
Adb21001101110	(	adb21001101110,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m011101_0	),
Adb21001101111	(	adb21001101111,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m011101_0	),
Adb21001110000	(	adb21001110000,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m011101_0	),
Adb21001110001	(	adb21001110001,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m011101_0	),
Adb21001110010	(	adb21001110010,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m011101_0	),
Adb21001110011	(	adb21001110011,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m011101_0	),
Adb21001110100	(	adb21001110100,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m011101_0	),
Adb21001110101	(	adb21001110101,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m011101_0	),
Adb21001110110	(	adb21001110110,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m011101_0	),
Adb21001110111	(	adb21001110111,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m011101_0	),
Adb21001111000	(	adb21001111000,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m011101_0	),
Adb21001111001	(	adb21001111001,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m011101_0	),
Adb21001111010	(	adb21001111010,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m011101_0	),
Adb21001111011	(	adb21001111011,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m011101_0	),
Adb21001111100	(	adb21001111100,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m011101_0	),
Adb21001111101	(	adb21001111101,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m011101_0	),
Adb21001111110	(	adb21001111110,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m011101_0	),
Adb21001111111	(	adb21001111111,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m011101_0	),
Adb21010000000	(	adb21010000000,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m010101_0	),
Adb21010000001	(	adb21010000001,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m010101_0	),
Adb21010000010	(	adb21010000010,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m010101_0	),
Adb21010000011	(	adb21010000011,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m010101_0	),
Adb21010000100	(	adb21010000100,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m010101_0	),
Adb21010000101	(	adb21010000101,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m010101_0	),
Adb21010000110	(	adb21010000110,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m010101_0	),
Adb21010000111	(	adb21010000111,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m010101_0	),
Adb21010001000	(	adb21010001000,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m010101_0	),
Adb21010001001	(	adb21010001001,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m010101_0	),
Adb21010001010	(	adb21010001010,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m010101_0	),
Adb21010001011	(	adb21010001011,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m010101_0	),
Adb21010001100	(	adb21010001100,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m010101_0	),
Adb21010001101	(	adb21010001101,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m010101_0	),
Adb21010001110	(	adb21010001110,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m010101_0	),
Adb21010001111	(	adb21010001111,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m010101_0	),
Adb21010010000	(	adb21010010000,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m010101_0	),
Adb21010010001	(	adb21010010001,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m010101_0	),
Adb21010010010	(	adb21010010010,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m010101_0	),
Adb21010010011	(	adb21010010011,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m010101_0	),
Adb21010010100	(	adb21010010100,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m010101_0	),
Adb21010010101	(	adb21010010101,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m010101_0	),
Adb21010010110	(	adb21010010110,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m010101_0	),
Adb21010010111	(	adb21010010111,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m010101_0	),
Adb21010011000	(	adb21010011000,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m010101_0	),
Adb21010011001	(	adb21010011001,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m010101_0	),
Adb21010011010	(	adb21010011010,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m010101_0	),
Adb21010011011	(	adb21010011011,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m010101_0	),
Adb21010011100	(	adb21010011100,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m010101_0	),
Adb21010011101	(	adb21010011101,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m010101_0	),
Adb21010011110	(	adb21010011110,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m010101_0	),
Adb21010011111	(	adb21010011111,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m010101_0	),
Adb21010100000	(	adb21010100000,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m010101_0	),
Adb21010100001	(	adb21010100001,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m010101_0	),
Adb21010100010	(	adb21010100010,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m010101_0	),
Adb21010100011	(	adb21010100011,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m010101_0	),
Adb21010100100	(	adb21010100100,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m010101_0	),
Adb21010100101	(	adb21010100101,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m010101_0	),
Adb21010100110	(	adb21010100110,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m010101_0	),
Adb21010100111	(	adb21010100111,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m010101_0	),
Adb21010101000	(	adb21010101000,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m010101_0	),
Adb21010101001	(	adb21010101001,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m010101_0	),
Adb21010101010	(	adb21010101010,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m010101_0	),
Adb21010101011	(	adb21010101011,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m010101_0	),
Adb21010101100	(	adb21010101100,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m010101_0	),
Adb21010101101	(	adb21010101101,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m010101_0	),
Adb21010101110	(	adb21010101110,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m010101_0	),
Adb21010101111	(	adb21010101111,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m010101_0	),
Adb21010110000	(	adb21010110000,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m010101_0	),
Adb21010110001	(	adb21010110001,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m010101_0	),
Adb21010110010	(	adb21010110010,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m010101_0	),
Adb21010110011	(	adb21010110011,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m010101_0	),
Adb21010110100	(	adb21010110100,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m010101_0	),
Adb21010110101	(	adb21010110101,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m010101_0	),
Adb21010110110	(	adb21010110110,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m010101_0	),
Adb21010110111	(	adb21010110111,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m010101_0	),
Adb21010111000	(	adb21010111000,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m010101_0	),
Adb21010111001	(	adb21010111001,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m010101_0	),
Adb21010111010	(	adb21010111010,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m010101_0	),
Adb21010111011	(	adb21010111011,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m010101_0	),
Adb21010111100	(	adb21010111100,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m010101_0	),
Adb21010111101	(	adb21010111101,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m010101_0	),
Adb21010111110	(	adb21010111110,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m010101_0	),
Adb21010111111	(	adb21010111111,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m010101_0	),
Adb21011000000	(	adb21011000000,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m010101_0	),
Adb21011000001	(	adb21011000001,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m010101_0	),
Adb21011000010	(	adb21011000010,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m010101_0	),
Adb21011000011	(	adb21011000011,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m010101_0	),
Adb21011000100	(	adb21011000100,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m010101_0	),
Adb21011000101	(	adb21011000101,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m010101_0	),
Adb21011000110	(	adb21011000110,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m010101_0	),
Adb21011000111	(	adb21011000111,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m010101_0	),
Adb21011001000	(	adb21011001000,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m010101_0	),
Adb21011001001	(	adb21011001001,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m010101_0	),
Adb21011001010	(	adb21011001010,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m010101_0	),
Adb21011001011	(	adb21011001011,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m010101_0	),
Adb21011001100	(	adb21011001100,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m010101_0	),
Adb21011001101	(	adb21011001101,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m010101_0	),
Adb21011001110	(	adb21011001110,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m010101_0	),
Adb21011001111	(	adb21011001111,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m010101_0	),
Adb21011010000	(	adb21011010000,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m010101_0	),
Adb21011010001	(	adb21011010001,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m010101_0	),
Adb21011010010	(	adb21011010010,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m010101_0	),
Adb21011010011	(	adb21011010011,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m010101_0	),
Adb21011010100	(	adb21011010100,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m010101_0	),
Adb21011010101	(	adb21011010101,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m010101_0	),
Adb21011010110	(	adb21011010110,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m010101_0	),
Adb21011010111	(	adb21011010111,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m010101_0	),
Adb21011011000	(	adb21011011000,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m010101_0	),
Adb21011011001	(	adb21011011001,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m010101_0	),
Adb21011011010	(	adb21011011010,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m010101_0	),
Adb21011011011	(	adb21011011011,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m010101_0	),
Adb21011011100	(	adb21011011100,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m010101_0	),
Adb21011011101	(	adb21011011101,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m010101_0	),
Adb21011011110	(	adb21011011110,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m010101_0	),
Adb21011011111	(	adb21011011111,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m010101_0	),
Adb21011100000	(	adb21011100000,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m010101_0	),
Adb21011100001	(	adb21011100001,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m010101_0	),
Adb21011100010	(	adb21011100010,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m010101_0	),
Adb21011100011	(	adb21011100011,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m010101_0	),
Adb21011100100	(	adb21011100100,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m010101_0	),
Adb21011100101	(	adb21011100101,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m010101_0	),
Adb21011100110	(	adb21011100110,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m010101_0	),
Adb21011100111	(	adb21011100111,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m010101_0	),
Adb21011101000	(	adb21011101000,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m010101_0	),
Adb21011101001	(	adb21011101001,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m010101_0	),
Adb21011101010	(	adb21011101010,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m010101_0	),
Adb21011101011	(	adb21011101011,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m010101_0	),
Adb21011101100	(	adb21011101100,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m010101_0	),
Adb21011101101	(	adb21011101101,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m010101_0	),
Adb21011101110	(	adb21011101110,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m010101_0	),
Adb21011101111	(	adb21011101111,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m010101_0	),
Adb21011110000	(	adb21011110000,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m010101_0	),
Adb21011110001	(	adb21011110001,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m010101_0	),
Adb21011110010	(	adb21011110010,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m010101_0	),
Adb21011110011	(	adb21011110011,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m010101_0	),
Adb21011110100	(	adb21011110100,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m010101_0	),
Adb21011110101	(	adb21011110101,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m010101_0	),
Adb21011110110	(	adb21011110110,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m010101_0	),
Adb21011110111	(	adb21011110111,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m010101_0	),
Adb21011111000	(	adb21011111000,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m010101_0	),
Adb21011111001	(	adb21011111001,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m010101_0	),
Adb21011111010	(	adb21011111010,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m010101_0	),
Adb21011111011	(	adb21011111011,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m010101_0	),
Adb21011111100	(	adb21011111100,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m010101_0	),
Adb21011111101	(	adb21011111101,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m010101_0	),
Adb21011111110	(	adb21011111110,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m010101_0	),
Adb21011111111	(	adb21011111111,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m010101_0	),
Adb21100000000	(	adb21100000000,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m001101_0	),
Adb21100000001	(	adb21100000001,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m001101_0	),
Adb21100000010	(	adb21100000010,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m001101_0	),
Adb21100000011	(	adb21100000011,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m001101_0	),
Adb21100000100	(	adb21100000100,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m001101_0	),
Adb21100000101	(	adb21100000101,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m001101_0	),
Adb21100000110	(	adb21100000110,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m001101_0	),
Adb21100000111	(	adb21100000111,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m001101_0	),
Adb21100001000	(	adb21100001000,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m001101_0	),
Adb21100001001	(	adb21100001001,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m001101_0	),
Adb21100001010	(	adb21100001010,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m001101_0	),
Adb21100001011	(	adb21100001011,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m001101_0	),
Adb21100001100	(	adb21100001100,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m001101_0	),
Adb21100001101	(	adb21100001101,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m001101_0	),
Adb21100001110	(	adb21100001110,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m001101_0	),
Adb21100001111	(	adb21100001111,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m001101_0	),
Adb21100010000	(	adb21100010000,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m001101_0	),
Adb21100010001	(	adb21100010001,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m001101_0	),
Adb21100010010	(	adb21100010010,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m001101_0	),
Adb21100010011	(	adb21100010011,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m001101_0	),
Adb21100010100	(	adb21100010100,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m001101_0	),
Adb21100010101	(	adb21100010101,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m001101_0	),
Adb21100010110	(	adb21100010110,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m001101_0	),
Adb21100010111	(	adb21100010111,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m001101_0	),
Adb21100011000	(	adb21100011000,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m001101_0	),
Adb21100011001	(	adb21100011001,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m001101_0	),
Adb21100011010	(	adb21100011010,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m001101_0	),
Adb21100011011	(	adb21100011011,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m001101_0	),
Adb21100011100	(	adb21100011100,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m001101_0	),
Adb21100011101	(	adb21100011101,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m001101_0	),
Adb21100011110	(	adb21100011110,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m001101_0	),
Adb21100011111	(	adb21100011111,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m001101_0	),
Adb21100100000	(	adb21100100000,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m001101_0	),
Adb21100100001	(	adb21100100001,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m001101_0	),
Adb21100100010	(	adb21100100010,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m001101_0	),
Adb21100100011	(	adb21100100011,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m001101_0	),
Adb21100100100	(	adb21100100100,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m001101_0	),
Adb21100100101	(	adb21100100101,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m001101_0	),
Adb21100100110	(	adb21100100110,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m001101_0	),
Adb21100100111	(	adb21100100111,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m001101_0	),
Adb21100101000	(	adb21100101000,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m001101_0	),
Adb21100101001	(	adb21100101001,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m001101_0	),
Adb21100101010	(	adb21100101010,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m001101_0	),
Adb21100101011	(	adb21100101011,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m001101_0	),
Adb21100101100	(	adb21100101100,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m001101_0	),
Adb21100101101	(	adb21100101101,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m001101_0	),
Adb21100101110	(	adb21100101110,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m001101_0	),
Adb21100101111	(	adb21100101111,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m001101_0	),
Adb21100110000	(	adb21100110000,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m001101_0	),
Adb21100110001	(	adb21100110001,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m001101_0	),
Adb21100110010	(	adb21100110010,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m001101_0	),
Adb21100110011	(	adb21100110011,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m001101_0	),
Adb21100110100	(	adb21100110100,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m001101_0	),
Adb21100110101	(	adb21100110101,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m001101_0	),
Adb21100110110	(	adb21100110110,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m001101_0	),
Adb21100110111	(	adb21100110111,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m001101_0	),
Adb21100111000	(	adb21100111000,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m001101_0	),
Adb21100111001	(	adb21100111001,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m001101_0	),
Adb21100111010	(	adb21100111010,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m001101_0	),
Adb21100111011	(	adb21100111011,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m001101_0	),
Adb21100111100	(	adb21100111100,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m001101_0	),
Adb21100111101	(	adb21100111101,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m001101_0	),
Adb21100111110	(	adb21100111110,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m001101_0	),
Adb21100111111	(	adb21100111111,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m001101_0	),
Adb21101000000	(	adb21101000000,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m001101_0	),
Adb21101000001	(	adb21101000001,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m001101_0	),
Adb21101000010	(	adb21101000010,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m001101_0	),
Adb21101000011	(	adb21101000011,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m001101_0	),
Adb21101000100	(	adb21101000100,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m001101_0	),
Adb21101000101	(	adb21101000101,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m001101_0	),
Adb21101000110	(	adb21101000110,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m001101_0	),
Adb21101000111	(	adb21101000111,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m001101_0	),
Adb21101001000	(	adb21101001000,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m001101_0	),
Adb21101001001	(	adb21101001001,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m001101_0	),
Adb21101001010	(	adb21101001010,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m001101_0	),
Adb21101001011	(	adb21101001011,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m001101_0	),
Adb21101001100	(	adb21101001100,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m001101_0	),
Adb21101001101	(	adb21101001101,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m001101_0	),
Adb21101001110	(	adb21101001110,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m001101_0	),
Adb21101001111	(	adb21101001111,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m001101_0	),
Adb21101010000	(	adb21101010000,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m001101_0	),
Adb21101010001	(	adb21101010001,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m001101_0	),
Adb21101010010	(	adb21101010010,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m001101_0	),
Adb21101010011	(	adb21101010011,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m001101_0	),
Adb21101010100	(	adb21101010100,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m001101_0	),
Adb21101010101	(	adb21101010101,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m001101_0	),
Adb21101010110	(	adb21101010110,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m001101_0	),
Adb21101010111	(	adb21101010111,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m001101_0	),
Adb21101011000	(	adb21101011000,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m001101_0	),
Adb21101011001	(	adb21101011001,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m001101_0	),
Adb21101011010	(	adb21101011010,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m001101_0	),
Adb21101011011	(	adb21101011011,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m001101_0	),
Adb21101011100	(	adb21101011100,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m001101_0	),
Adb21101011101	(	adb21101011101,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m001101_0	),
Adb21101011110	(	adb21101011110,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m001101_0	),
Adb21101011111	(	adb21101011111,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m001101_0	),
Adb21101100000	(	adb21101100000,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m001101_0	),
Adb21101100001	(	adb21101100001,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m001101_0	),
Adb21101100010	(	adb21101100010,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m001101_0	),
Adb21101100011	(	adb21101100011,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m001101_0	),
Adb21101100100	(	adb21101100100,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m001101_0	),
Adb21101100101	(	adb21101100101,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m001101_0	),
Adb21101100110	(	adb21101100110,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m001101_0	),
Adb21101100111	(	adb21101100111,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m001101_0	),
Adb21101101000	(	adb21101101000,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m001101_0	),
Adb21101101001	(	adb21101101001,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m001101_0	),
Adb21101101010	(	adb21101101010,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m001101_0	),
Adb21101101011	(	adb21101101011,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m001101_0	),
Adb21101101100	(	adb21101101100,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m001101_0	),
Adb21101101101	(	adb21101101101,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m001101_0	),
Adb21101101110	(	adb21101101110,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m001101_0	),
Adb21101101111	(	adb21101101111,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m001101_0	),
Adb21101110000	(	adb21101110000,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m001101_0	),
Adb21101110001	(	adb21101110001,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m001101_0	),
Adb21101110010	(	adb21101110010,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m001101_0	),
Adb21101110011	(	adb21101110011,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m001101_0	),
Adb21101110100	(	adb21101110100,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m001101_0	),
Adb21101110101	(	adb21101110101,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m001101_0	),
Adb21101110110	(	adb21101110110,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m001101_0	),
Adb21101110111	(	adb21101110111,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m001101_0	),
Adb21101111000	(	adb21101111000,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m001101_0	),
Adb21101111001	(	adb21101111001,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m001101_0	),
Adb21101111010	(	adb21101111010,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m001101_0	),
Adb21101111011	(	adb21101111011,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m001101_0	),
Adb21101111100	(	adb21101111100,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m001101_0	),
Adb21101111101	(	adb21101111101,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m001101_0	),
Adb21101111110	(	adb21101111110,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m001101_0	),
Adb21101111111	(	adb21101111111,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m001101_0	),
Adb21110000000	(	adb21110000000,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m000101_0	),
Adb21110000001	(	adb21110000001,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m000101_0	),
Adb21110000010	(	adb21110000010,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m000101_0	),
Adb21110000011	(	adb21110000011,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m000101_0	),
Adb21110000100	(	adb21110000100,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m000101_0	),
Adb21110000101	(	adb21110000101,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m000101_0	),
Adb21110000110	(	adb21110000110,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m000101_0	),
Adb21110000111	(	adb21110000111,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m000101_0	),
Adb21110001000	(	adb21110001000,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m000101_0	),
Adb21110001001	(	adb21110001001,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m000101_0	),
Adb21110001010	(	adb21110001010,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m000101_0	),
Adb21110001011	(	adb21110001011,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m000101_0	),
Adb21110001100	(	adb21110001100,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m000101_0	),
Adb21110001101	(	adb21110001101,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m000101_0	),
Adb21110001110	(	adb21110001110,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m000101_0	),
Adb21110001111	(	adb21110001111,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m000101_0	),
Adb21110010000	(	adb21110010000,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m000101_0	),
Adb21110010001	(	adb21110010001,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m000101_0	),
Adb21110010010	(	adb21110010010,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m000101_0	),
Adb21110010011	(	adb21110010011,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m000101_0	),
Adb21110010100	(	adb21110010100,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m000101_0	),
Adb21110010101	(	adb21110010101,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m000101_0	),
Adb21110010110	(	adb21110010110,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m000101_0	),
Adb21110010111	(	adb21110010111,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m000101_0	),
Adb21110011000	(	adb21110011000,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m000101_0	),
Adb21110011001	(	adb21110011001,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m000101_0	),
Adb21110011010	(	adb21110011010,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m000101_0	),
Adb21110011011	(	adb21110011011,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m000101_0	),
Adb21110011100	(	adb21110011100,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m000101_0	),
Adb21110011101	(	adb21110011101,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m000101_0	),
Adb21110011110	(	adb21110011110,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m000101_0	),
Adb21110011111	(	adb21110011111,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m000101_0	),
Adb21110100000	(	adb21110100000,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m000101_0	),
Adb21110100001	(	adb21110100001,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m000101_0	),
Adb21110100010	(	adb21110100010,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m000101_0	),
Adb21110100011	(	adb21110100011,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m000101_0	),
Adb21110100100	(	adb21110100100,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m000101_0	),
Adb21110100101	(	adb21110100101,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m000101_0	),
Adb21110100110	(	adb21110100110,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m000101_0	),
Adb21110100111	(	adb21110100111,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m000101_0	),
Adb21110101000	(	adb21110101000,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m000101_0	),
Adb21110101001	(	adb21110101001,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m000101_0	),
Adb21110101010	(	adb21110101010,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m000101_0	),
Adb21110101011	(	adb21110101011,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m000101_0	),
Adb21110101100	(	adb21110101100,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m000101_0	),
Adb21110101101	(	adb21110101101,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m000101_0	),
Adb21110101110	(	adb21110101110,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m000101_0	),
Adb21110101111	(	adb21110101111,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m000101_0	),
Adb21110110000	(	adb21110110000,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m000101_0	),
Adb21110110001	(	adb21110110001,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m000101_0	),
Adb21110110010	(	adb21110110010,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m000101_0	),
Adb21110110011	(	adb21110110011,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m000101_0	),
Adb21110110100	(	adb21110110100,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m000101_0	),
Adb21110110101	(	adb21110110101,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m000101_0	),
Adb21110110110	(	adb21110110110,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m000101_0	),
Adb21110110111	(	adb21110110111,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m000101_0	),
Adb21110111000	(	adb21110111000,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m000101_0	),
Adb21110111001	(	adb21110111001,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m000101_0	),
Adb21110111010	(	adb21110111010,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m000101_0	),
Adb21110111011	(	adb21110111011,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m000101_0	),
Adb21110111100	(	adb21110111100,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m000101_0	),
Adb21110111101	(	adb21110111101,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m000101_0	),
Adb21110111110	(	adb21110111110,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m000101_0	),
Adb21110111111	(	adb21110111111,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m000101_0	),
Adb21111000000	(	adb21111000000,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m000101_0	),
Adb21111000001	(	adb21111000001,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m000101_0	),
Adb21111000010	(	adb21111000010,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m000101_0	),
Adb21111000011	(	adb21111000011,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m000101_0	),
Adb21111000100	(	adb21111000100,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m000101_0	),
Adb21111000101	(	adb21111000101,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m000101_0	),
Adb21111000110	(	adb21111000110,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m000101_0	),
Adb21111000111	(	adb21111000111,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m000101_0	),
Adb21111001000	(	adb21111001000,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m000101_0	),
Adb21111001001	(	adb21111001001,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m000101_0	),
Adb21111001010	(	adb21111001010,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m000101_0	),
Adb21111001011	(	adb21111001011,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m000101_0	),
Adb21111001100	(	adb21111001100,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m000101_0	),
Adb21111001101	(	adb21111001101,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m000101_0	),
Adb21111001110	(	adb21111001110,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m000101_0	),
Adb21111001111	(	adb21111001111,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m000101_0	),
Adb21111010000	(	adb21111010000,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m000101_0	),
Adb21111010001	(	adb21111010001,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m000101_0	),
Adb21111010010	(	adb21111010010,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m000101_0	),
Adb21111010011	(	adb21111010011,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m000101_0	),
Adb21111010100	(	adb21111010100,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m000101_0	),
Adb21111010101	(	adb21111010101,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m000101_0	),
Adb21111010110	(	adb21111010110,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m000101_0	),
Adb21111010111	(	adb21111010111,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m000101_0	),
Adb21111011000	(	adb21111011000,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m000101_0	),
Adb21111011001	(	adb21111011001,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m000101_0	),
Adb21111011010	(	adb21111011010,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m000101_0	),
Adb21111011011	(	adb21111011011,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m000101_0	),
Adb21111011100	(	adb21111011100,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m000101_0	),
Adb21111011101	(	adb21111011101,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m000101_0	),
Adb21111011110	(	adb21111011110,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m000101_0	),
Adb21111011111	(	adb21111011111,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m000101_0	),
Adb21111100000	(	adb21111100000,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m000101_0	),
Adb21111100001	(	adb21111100001,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m000101_0	),
Adb21111100010	(	adb21111100010,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m000101_0	),
Adb21111100011	(	adb21111100011,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m000101_0	),
Adb21111100100	(	adb21111100100,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m000101_0	),
Adb21111100101	(	adb21111100101,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m000101_0	),
Adb21111100110	(	adb21111100110,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m000101_0	),
Adb21111100111	(	adb21111100111,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m000101_0	),
Adb21111101000	(	adb21111101000,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m000101_0	),
Adb21111101001	(	adb21111101001,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m000101_0	),
Adb21111101010	(	adb21111101010,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m000101_0	),
Adb21111101011	(	adb21111101011,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m000101_0	),
Adb21111101100	(	adb21111101100,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m000101_0	),
Adb21111101101	(	adb21111101101,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m000101_0	),
Adb21111101110	(	adb21111101110,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m000101_0	),
Adb21111101111	(	adb21111101111,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m000101_0	),
Adb21111110000	(	adb21111110000,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m000101_0	),
Adb21111110001	(	adb21111110001,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m000101_0	),
Adb21111110010	(	adb21111110010,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m000101_0	),
Adb21111110011	(	adb21111110011,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m000101_0	),
Adb21111110100	(	adb21111110100,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m000101_0	),
Adb21111110101	(	adb21111110101,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m000101_0	),
Adb21111110110	(	adb21111110110,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m000101_0	),
Adb21111110111	(	adb21111110111,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m000101_0	),
Adb21111111000	(	adb21111111000,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m000101_0	),
Adb21111111001	(	adb21111111001,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m000101_0	),
Adb21111111010	(	adb21111111010,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m000101_0	),
Adb21111111011	(	adb21111111011,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m000101_0	),
Adb21111111100	(	adb21111111100,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m000101_0	),
Adb21111111101	(	adb21111111101,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m000101_0	),
Adb21111111110	(	adb21111111110,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m000101_0	),
Adb21111111111	(	adb21111111111,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m000101_0	),
       Adb300(adb300,n0011,n0010,n0009,dbv1),
       Adb301(adb301,n0011,n0010,m0009,m0013),
       Adb310(adb310,n0011,m0010,n0009,dbv1),
       Adb311(adb311,n0011,m0010,m0009,dbv0),
Adb30000000000	(	adb30000000000,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m111100_0	),
Adb30000000001	(	adb30000000001,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m111100_0	),
Adb30000000010	(	adb30000000010,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m111100_0	),
Adb30000000011	(	adb30000000011,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m111100_0	),
Adb30000000100	(	adb30000000100,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m111100_0	),
Adb30000000101	(	adb30000000101,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m111100_0	),
Adb30000000110	(	adb30000000110,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m111100_0	),
Adb30000000111	(	adb30000000111,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m111100_0	),
Adb30000001000	(	adb30000001000,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m111100_0	),
Adb30000001001	(	adb30000001001,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m111100_0	),
Adb30000001010	(	adb30000001010,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m111100_0	),
Adb30000001011	(	adb30000001011,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m111100_0	),
Adb30000001100	(	adb30000001100,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m111100_0	),
Adb30000001101	(	adb30000001101,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m111100_0	),
Adb30000001110	(	adb30000001110,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m111100_0	),
Adb30000001111	(	adb30000001111,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m111100_0	),
Adb30000010000	(	adb30000010000,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m111100_0	),
Adb30000010001	(	adb30000010001,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m111100_0	),
Adb30000010010	(	adb30000010010,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m111100_0	),
Adb30000010011	(	adb30000010011,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m111100_0	),
Adb30000010100	(	adb30000010100,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m111100_0	),
Adb30000010101	(	adb30000010101,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m111100_0	),
Adb30000010110	(	adb30000010110,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m111100_0	),
Adb30000010111	(	adb30000010111,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m111100_0	),
Adb30000011000	(	adb30000011000,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m111100_0	),
Adb30000011001	(	adb30000011001,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m111100_0	),
Adb30000011010	(	adb30000011010,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m111100_0	),
Adb30000011011	(	adb30000011011,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m111100_0	),
Adb30000011100	(	adb30000011100,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m111100_0	),
Adb30000011101	(	adb30000011101,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m111100_0	),
Adb30000011110	(	adb30000011110,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m111100_0	),
Adb30000011111	(	adb30000011111,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m111100_0	),
Adb30000100000	(	adb30000100000,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m111100_0	),
Adb30000100001	(	adb30000100001,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m111100_0	),
Adb30000100010	(	adb30000100010,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m111100_0	),
Adb30000100011	(	adb30000100011,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m111100_0	),
Adb30000100100	(	adb30000100100,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m111100_0	),
Adb30000100101	(	adb30000100101,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m111100_0	),
Adb30000100110	(	adb30000100110,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m111100_0	),
Adb30000100111	(	adb30000100111,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m111100_0	),
Adb30000101000	(	adb30000101000,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m111100_0	),
Adb30000101001	(	adb30000101001,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m111100_0	),
Adb30000101010	(	adb30000101010,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m111100_0	),
Adb30000101011	(	adb30000101011,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m111100_0	),
Adb30000101100	(	adb30000101100,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m111100_0	),
Adb30000101101	(	adb30000101101,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m111100_0	),
Adb30000101110	(	adb30000101110,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m111100_0	),
Adb30000101111	(	adb30000101111,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m111100_0	),
Adb30000110000	(	adb30000110000,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m111100_0	),
Adb30000110001	(	adb30000110001,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m111100_0	),
Adb30000110010	(	adb30000110010,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m111100_0	),
Adb30000110011	(	adb30000110011,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m111100_0	),
Adb30000110100	(	adb30000110100,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m111100_0	),
Adb30000110101	(	adb30000110101,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m111100_0	),
Adb30000110110	(	adb30000110110,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m111100_0	),
Adb30000110111	(	adb30000110111,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m111100_0	),
Adb30000111000	(	adb30000111000,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m111100_0	),
Adb30000111001	(	adb30000111001,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m111100_0	),
Adb30000111010	(	adb30000111010,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m111100_0	),
Adb30000111011	(	adb30000111011,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m111100_0	),
Adb30000111100	(	adb30000111100,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m111100_0	),
Adb30000111101	(	adb30000111101,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m111100_0	),
Adb30000111110	(	adb30000111110,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m111100_0	),
Adb30000111111	(	adb30000111111,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m111100_0	),
Adb30001000000	(	adb30001000000,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m111100_0	),
Adb30001000001	(	adb30001000001,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m111100_0	),
Adb30001000010	(	adb30001000010,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m111100_0	),
Adb30001000011	(	adb30001000011,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m111100_0	),
Adb30001000100	(	adb30001000100,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m111100_0	),
Adb30001000101	(	adb30001000101,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m111100_0	),
Adb30001000110	(	adb30001000110,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m111100_0	),
Adb30001000111	(	adb30001000111,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m111100_0	),
Adb30001001000	(	adb30001001000,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m111100_0	),
Adb30001001001	(	adb30001001001,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m111100_0	),
Adb30001001010	(	adb30001001010,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m111100_0	),
Adb30001001011	(	adb30001001011,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m111100_0	),
Adb30001001100	(	adb30001001100,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m111100_0	),
Adb30001001101	(	adb30001001101,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m111100_0	),
Adb30001001110	(	adb30001001110,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m111100_0	),
Adb30001001111	(	adb30001001111,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m111100_0	),
Adb30001010000	(	adb30001010000,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m111100_0	),
Adb30001010001	(	adb30001010001,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m111100_0	),
Adb30001010010	(	adb30001010010,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m111100_0	),
Adb30001010011	(	adb30001010011,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m111100_0	),
Adb30001010100	(	adb30001010100,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m111100_0	),
Adb30001010101	(	adb30001010101,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m111100_0	),
Adb30001010110	(	adb30001010110,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m111100_0	),
Adb30001010111	(	adb30001010111,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m111100_0	),
Adb30001011000	(	adb30001011000,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m111100_0	),
Adb30001011001	(	adb30001011001,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m111100_0	),
Adb30001011010	(	adb30001011010,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m111100_0	),
Adb30001011011	(	adb30001011011,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m111100_0	),
Adb30001011100	(	adb30001011100,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m111100_0	),
Adb30001011101	(	adb30001011101,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m111100_0	),
Adb30001011110	(	adb30001011110,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m111100_0	),
Adb30001011111	(	adb30001011111,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m111100_0	),
Adb30001100000	(	adb30001100000,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m111100_0	),
Adb30001100001	(	adb30001100001,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m111100_0	),
Adb30001100010	(	adb30001100010,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m111100_0	),
Adb30001100011	(	adb30001100011,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m111100_0	),
Adb30001100100	(	adb30001100100,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m111100_0	),
Adb30001100101	(	adb30001100101,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m111100_0	),
Adb30001100110	(	adb30001100110,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m111100_0	),
Adb30001100111	(	adb30001100111,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m111100_0	),
Adb30001101000	(	adb30001101000,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m111100_0	),
Adb30001101001	(	adb30001101001,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m111100_0	),
Adb30001101010	(	adb30001101010,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m111100_0	),
Adb30001101011	(	adb30001101011,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m111100_0	),
Adb30001101100	(	adb30001101100,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m111100_0	),
Adb30001101101	(	adb30001101101,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m111100_0	),
Adb30001101110	(	adb30001101110,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m111100_0	),
Adb30001101111	(	adb30001101111,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m111100_0	),
Adb30001110000	(	adb30001110000,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m111100_0	),
Adb30001110001	(	adb30001110001,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m111100_0	),
Adb30001110010	(	adb30001110010,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m111100_0	),
Adb30001110011	(	adb30001110011,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m111100_0	),
Adb30001110100	(	adb30001110100,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m111100_0	),
Adb30001110101	(	adb30001110101,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m111100_0	),
Adb30001110110	(	adb30001110110,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m111100_0	),
Adb30001110111	(	adb30001110111,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m111100_0	),
Adb30001111000	(	adb30001111000,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m111100_0	),
Adb30001111001	(	adb30001111001,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m111100_0	),
Adb30001111010	(	adb30001111010,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m111100_0	),
Adb30001111011	(	adb30001111011,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m111100_0	),
Adb30001111100	(	adb30001111100,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m111100_0	),
Adb30001111101	(	adb30001111101,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m111100_0	),
Adb30001111110	(	adb30001111110,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m111100_0	),
Adb30001111111	(	adb30001111111,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m111100_0	),
Adb30010000000	(	adb30010000000,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m110100_0	),
Adb30010000001	(	adb30010000001,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m110100_0	),
Adb30010000010	(	adb30010000010,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m110100_0	),
Adb30010000011	(	adb30010000011,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m110100_0	),
Adb30010000100	(	adb30010000100,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m110100_0	),
Adb30010000101	(	adb30010000101,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m110100_0	),
Adb30010000110	(	adb30010000110,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m110100_0	),
Adb30010000111	(	adb30010000111,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m110100_0	),
Adb30010001000	(	adb30010001000,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m110100_0	),
Adb30010001001	(	adb30010001001,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m110100_0	),
Adb30010001010	(	adb30010001010,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m110100_0	),
Adb30010001011	(	adb30010001011,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m110100_0	),
Adb30010001100	(	adb30010001100,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m110100_0	),
Adb30010001101	(	adb30010001101,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m110100_0	),
Adb30010001110	(	adb30010001110,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m110100_0	),
Adb30010001111	(	adb30010001111,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m110100_0	),
Adb30010010000	(	adb30010010000,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m110100_0	),
Adb30010010001	(	adb30010010001,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m110100_0	),
Adb30010010010	(	adb30010010010,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m110100_0	),
Adb30010010011	(	adb30010010011,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m110100_0	),
Adb30010010100	(	adb30010010100,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m110100_0	),
Adb30010010101	(	adb30010010101,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m110100_0	),
Adb30010010110	(	adb30010010110,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m110100_0	),
Adb30010010111	(	adb30010010111,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m110100_0	),
Adb30010011000	(	adb30010011000,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m110100_0	),
Adb30010011001	(	adb30010011001,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m110100_0	),
Adb30010011010	(	adb30010011010,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m110100_0	),
Adb30010011011	(	adb30010011011,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m110100_0	),
Adb30010011100	(	adb30010011100,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m110100_0	),
Adb30010011101	(	adb30010011101,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m110100_0	),
Adb30010011110	(	adb30010011110,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m110100_0	),
Adb30010011111	(	adb30010011111,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m110100_0	),
Adb30010100000	(	adb30010100000,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m110100_0	),
Adb30010100001	(	adb30010100001,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m110100_0	),
Adb30010100010	(	adb30010100010,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m110100_0	),
Adb30010100011	(	adb30010100011,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m110100_0	),
Adb30010100100	(	adb30010100100,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m110100_0	),
Adb30010100101	(	adb30010100101,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m110100_0	),
Adb30010100110	(	adb30010100110,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m110100_0	),
Adb30010100111	(	adb30010100111,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m110100_0	),
Adb30010101000	(	adb30010101000,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m110100_0	),
Adb30010101001	(	adb30010101001,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m110100_0	),
Adb30010101010	(	adb30010101010,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m110100_0	),
Adb30010101011	(	adb30010101011,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m110100_0	),
Adb30010101100	(	adb30010101100,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m110100_0	),
Adb30010101101	(	adb30010101101,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m110100_0	),
Adb30010101110	(	adb30010101110,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m110100_0	),
Adb30010101111	(	adb30010101111,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m110100_0	),
Adb30010110000	(	adb30010110000,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m110100_0	),
Adb30010110001	(	adb30010110001,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m110100_0	),
Adb30010110010	(	adb30010110010,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m110100_0	),
Adb30010110011	(	adb30010110011,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m110100_0	),
Adb30010110100	(	adb30010110100,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m110100_0	),
Adb30010110101	(	adb30010110101,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m110100_0	),
Adb30010110110	(	adb30010110110,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m110100_0	),
Adb30010110111	(	adb30010110111,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m110100_0	),
Adb30010111000	(	adb30010111000,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m110100_0	),
Adb30010111001	(	adb30010111001,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m110100_0	),
Adb30010111010	(	adb30010111010,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m110100_0	),
Adb30010111011	(	adb30010111011,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m110100_0	),
Adb30010111100	(	adb30010111100,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m110100_0	),
Adb30010111101	(	adb30010111101,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m110100_0	),
Adb30010111110	(	adb30010111110,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m110100_0	),
Adb30010111111	(	adb30010111111,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m110100_0	),
Adb30011000000	(	adb30011000000,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m110100_0	),
Adb30011000001	(	adb30011000001,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m110100_0	),
Adb30011000010	(	adb30011000010,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m110100_0	),
Adb30011000011	(	adb30011000011,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m110100_0	),
Adb30011000100	(	adb30011000100,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m110100_0	),
Adb30011000101	(	adb30011000101,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m110100_0	),
Adb30011000110	(	adb30011000110,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m110100_0	),
Adb30011000111	(	adb30011000111,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m110100_0	),
Adb30011001000	(	adb30011001000,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m110100_0	),
Adb30011001001	(	adb30011001001,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m110100_0	),
Adb30011001010	(	adb30011001010,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m110100_0	),
Adb30011001011	(	adb30011001011,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m110100_0	),
Adb30011001100	(	adb30011001100,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m110100_0	),
Adb30011001101	(	adb30011001101,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m110100_0	),
Adb30011001110	(	adb30011001110,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m110100_0	),
Adb30011001111	(	adb30011001111,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m110100_0	),
Adb30011010000	(	adb30011010000,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m110100_0	),
Adb30011010001	(	adb30011010001,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m110100_0	),
Adb30011010010	(	adb30011010010,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m110100_0	),
Adb30011010011	(	adb30011010011,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m110100_0	),
Adb30011010100	(	adb30011010100,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m110100_0	),
Adb30011010101	(	adb30011010101,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m110100_0	),
Adb30011010110	(	adb30011010110,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m110100_0	),
Adb30011010111	(	adb30011010111,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m110100_0	),
Adb30011011000	(	adb30011011000,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m110100_0	),
Adb30011011001	(	adb30011011001,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m110100_0	),
Adb30011011010	(	adb30011011010,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m110100_0	),
Adb30011011011	(	adb30011011011,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m110100_0	),
Adb30011011100	(	adb30011011100,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m110100_0	),
Adb30011011101	(	adb30011011101,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m110100_0	),
Adb30011011110	(	adb30011011110,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m110100_0	),
Adb30011011111	(	adb30011011111,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m110100_0	),
Adb30011100000	(	adb30011100000,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m110100_0	),
Adb30011100001	(	adb30011100001,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m110100_0	),
Adb30011100010	(	adb30011100010,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m110100_0	),
Adb30011100011	(	adb30011100011,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m110100_0	),
Adb30011100100	(	adb30011100100,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m110100_0	),
Adb30011100101	(	adb30011100101,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m110100_0	),
Adb30011100110	(	adb30011100110,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m110100_0	),
Adb30011100111	(	adb30011100111,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m110100_0	),
Adb30011101000	(	adb30011101000,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m110100_0	),
Adb30011101001	(	adb30011101001,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m110100_0	),
Adb30011101010	(	adb30011101010,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m110100_0	),
Adb30011101011	(	adb30011101011,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m110100_0	),
Adb30011101100	(	adb30011101100,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m110100_0	),
Adb30011101101	(	adb30011101101,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m110100_0	),
Adb30011101110	(	adb30011101110,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m110100_0	),
Adb30011101111	(	adb30011101111,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m110100_0	),
Adb30011110000	(	adb30011110000,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m110100_0	),
Adb30011110001	(	adb30011110001,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m110100_0	),
Adb30011110010	(	adb30011110010,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m110100_0	),
Adb30011110011	(	adb30011110011,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m110100_0	),
Adb30011110100	(	adb30011110100,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m110100_0	),
Adb30011110101	(	adb30011110101,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m110100_0	),
Adb30011110110	(	adb30011110110,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m110100_0	),
Adb30011110111	(	adb30011110111,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m110100_0	),
Adb30011111000	(	adb30011111000,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m110100_0	),
Adb30011111001	(	adb30011111001,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m110100_0	),
Adb30011111010	(	adb30011111010,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m110100_0	),
Adb30011111011	(	adb30011111011,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m110100_0	),
Adb30011111100	(	adb30011111100,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m110100_0	),
Adb30011111101	(	adb30011111101,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m110100_0	),
Adb30011111110	(	adb30011111110,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m110100_0	),
Adb30011111111	(	adb30011111111,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m110100_0	),
Adb30100000000	(	adb30100000000,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m101100_0	),
Adb30100000001	(	adb30100000001,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m101100_0	),
Adb30100000010	(	adb30100000010,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m101100_0	),
Adb30100000011	(	adb30100000011,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m101100_0	),
Adb30100000100	(	adb30100000100,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m101100_0	),
Adb30100000101	(	adb30100000101,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m101100_0	),
Adb30100000110	(	adb30100000110,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m101100_0	),
Adb30100000111	(	adb30100000111,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m101100_0	),
Adb30100001000	(	adb30100001000,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m101100_0	),
Adb30100001001	(	adb30100001001,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m101100_0	),
Adb30100001010	(	adb30100001010,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m101100_0	),
Adb30100001011	(	adb30100001011,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m101100_0	),
Adb30100001100	(	adb30100001100,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m101100_0	),
Adb30100001101	(	adb30100001101,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m101100_0	),
Adb30100001110	(	adb30100001110,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m101100_0	),
Adb30100001111	(	adb30100001111,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m101100_0	),
Adb30100010000	(	adb30100010000,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m101100_0	),
Adb30100010001	(	adb30100010001,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m101100_0	),
Adb30100010010	(	adb30100010010,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m101100_0	),
Adb30100010011	(	adb30100010011,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m101100_0	),
Adb30100010100	(	adb30100010100,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m101100_0	),
Adb30100010101	(	adb30100010101,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m101100_0	),
Adb30100010110	(	adb30100010110,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m101100_0	),
Adb30100010111	(	adb30100010111,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m101100_0	),
Adb30100011000	(	adb30100011000,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m101100_0	),
Adb30100011001	(	adb30100011001,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m101100_0	),
Adb30100011010	(	adb30100011010,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m101100_0	),
Adb30100011011	(	adb30100011011,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m101100_0	),
Adb30100011100	(	adb30100011100,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m101100_0	),
Adb30100011101	(	adb30100011101,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m101100_0	),
Adb30100011110	(	adb30100011110,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m101100_0	),
Adb30100011111	(	adb30100011111,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m101100_0	),
Adb30100100000	(	adb30100100000,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m101100_0	),
Adb30100100001	(	adb30100100001,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m101100_0	),
Adb30100100010	(	adb30100100010,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m101100_0	),
Adb30100100011	(	adb30100100011,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m101100_0	),
Adb30100100100	(	adb30100100100,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m101100_0	),
Adb30100100101	(	adb30100100101,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m101100_0	),
Adb30100100110	(	adb30100100110,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m101100_0	),
Adb30100100111	(	adb30100100111,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m101100_0	),
Adb30100101000	(	adb30100101000,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m101100_0	),
Adb30100101001	(	adb30100101001,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m101100_0	),
Adb30100101010	(	adb30100101010,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m101100_0	),
Adb30100101011	(	adb30100101011,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m101100_0	),
Adb30100101100	(	adb30100101100,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m101100_0	),
Adb30100101101	(	adb30100101101,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m101100_0	),
Adb30100101110	(	adb30100101110,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m101100_0	),
Adb30100101111	(	adb30100101111,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m101100_0	),
Adb30100110000	(	adb30100110000,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m101100_0	),
Adb30100110001	(	adb30100110001,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m101100_0	),
Adb30100110010	(	adb30100110010,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m101100_0	),
Adb30100110011	(	adb30100110011,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m101100_0	),
Adb30100110100	(	adb30100110100,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m101100_0	),
Adb30100110101	(	adb30100110101,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m101100_0	),
Adb30100110110	(	adb30100110110,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m101100_0	),
Adb30100110111	(	adb30100110111,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m101100_0	),
Adb30100111000	(	adb30100111000,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m101100_0	),
Adb30100111001	(	adb30100111001,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m101100_0	),
Adb30100111010	(	adb30100111010,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m101100_0	),
Adb30100111011	(	adb30100111011,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m101100_0	),
Adb30100111100	(	adb30100111100,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m101100_0	),
Adb30100111101	(	adb30100111101,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m101100_0	),
Adb30100111110	(	adb30100111110,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m101100_0	),
Adb30100111111	(	adb30100111111,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m101100_0	),
Adb30101000000	(	adb30101000000,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m101100_0	),
Adb30101000001	(	adb30101000001,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m101100_0	),
Adb30101000010	(	adb30101000010,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m101100_0	),
Adb30101000011	(	adb30101000011,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m101100_0	),
Adb30101000100	(	adb30101000100,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m101100_0	),
Adb30101000101	(	adb30101000101,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m101100_0	),
Adb30101000110	(	adb30101000110,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m101100_0	),
Adb30101000111	(	adb30101000111,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m101100_0	),
Adb30101001000	(	adb30101001000,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m101100_0	),
Adb30101001001	(	adb30101001001,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m101100_0	),
Adb30101001010	(	adb30101001010,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m101100_0	),
Adb30101001011	(	adb30101001011,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m101100_0	),
Adb30101001100	(	adb30101001100,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m101100_0	),
Adb30101001101	(	adb30101001101,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m101100_0	),
Adb30101001110	(	adb30101001110,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m101100_0	),
Adb30101001111	(	adb30101001111,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m101100_0	),
Adb30101010000	(	adb30101010000,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m101100_0	),
Adb30101010001	(	adb30101010001,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m101100_0	),
Adb30101010010	(	adb30101010010,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m101100_0	),
Adb30101010011	(	adb30101010011,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m101100_0	),
Adb30101010100	(	adb30101010100,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m101100_0	),
Adb30101010101	(	adb30101010101,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m101100_0	),
Adb30101010110	(	adb30101010110,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m101100_0	),
Adb30101010111	(	adb30101010111,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m101100_0	),
Adb30101011000	(	adb30101011000,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m101100_0	),
Adb30101011001	(	adb30101011001,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m101100_0	),
Adb30101011010	(	adb30101011010,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m101100_0	),
Adb30101011011	(	adb30101011011,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m101100_0	),
Adb30101011100	(	adb30101011100,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m101100_0	),
Adb30101011101	(	adb30101011101,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m101100_0	),
Adb30101011110	(	adb30101011110,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m101100_0	),
Adb30101011111	(	adb30101011111,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m101100_0	),
Adb30101100000	(	adb30101100000,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m101100_0	),
Adb30101100001	(	adb30101100001,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m101100_0	),
Adb30101100010	(	adb30101100010,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m101100_0	),
Adb30101100011	(	adb30101100011,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m101100_0	),
Adb30101100100	(	adb30101100100,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m101100_0	),
Adb30101100101	(	adb30101100101,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m101100_0	),
Adb30101100110	(	adb30101100110,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m101100_0	),
Adb30101100111	(	adb30101100111,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m101100_0	),
Adb30101101000	(	adb30101101000,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m101100_0	),
Adb30101101001	(	adb30101101001,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m101100_0	),
Adb30101101010	(	adb30101101010,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m101100_0	),
Adb30101101011	(	adb30101101011,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m101100_0	),
Adb30101101100	(	adb30101101100,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m101100_0	),
Adb30101101101	(	adb30101101101,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m101100_0	),
Adb30101101110	(	adb30101101110,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m101100_0	),
Adb30101101111	(	adb30101101111,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m101100_0	),
Adb30101110000	(	adb30101110000,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m101100_0	),
Adb30101110001	(	adb30101110001,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m101100_0	),
Adb30101110010	(	adb30101110010,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m101100_0	),
Adb30101110011	(	adb30101110011,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m101100_0	),
Adb30101110100	(	adb30101110100,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m101100_0	),
Adb30101110101	(	adb30101110101,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m101100_0	),
Adb30101110110	(	adb30101110110,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m101100_0	),
Adb30101110111	(	adb30101110111,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m101100_0	),
Adb30101111000	(	adb30101111000,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m101100_0	),
Adb30101111001	(	adb30101111001,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m101100_0	),
Adb30101111010	(	adb30101111010,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m101100_0	),
Adb30101111011	(	adb30101111011,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m101100_0	),
Adb30101111100	(	adb30101111100,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m101100_0	),
Adb30101111101	(	adb30101111101,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m101100_0	),
Adb30101111110	(	adb30101111110,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m101100_0	),
Adb30101111111	(	adb30101111111,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m101100_0	),
Adb30110000000	(	adb30110000000,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m100100_0	),
Adb30110000001	(	adb30110000001,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m100100_0	),
Adb30110000010	(	adb30110000010,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m100100_0	),
Adb30110000011	(	adb30110000011,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m100100_0	),
Adb30110000100	(	adb30110000100,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m100100_0	),
Adb30110000101	(	adb30110000101,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m100100_0	),
Adb30110000110	(	adb30110000110,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m100100_0	),
Adb30110000111	(	adb30110000111,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m100100_0	),
Adb30110001000	(	adb30110001000,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m100100_0	),
Adb30110001001	(	adb30110001001,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m100100_0	),
Adb30110001010	(	adb30110001010,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m100100_0	),
Adb30110001011	(	adb30110001011,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m100100_0	),
Adb30110001100	(	adb30110001100,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m100100_0	),
Adb30110001101	(	adb30110001101,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m100100_0	),
Adb30110001110	(	adb30110001110,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m100100_0	),
Adb30110001111	(	adb30110001111,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m100100_0	),
Adb30110010000	(	adb30110010000,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m100100_0	),
Adb30110010001	(	adb30110010001,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m100100_0	),
Adb30110010010	(	adb30110010010,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m100100_0	),
Adb30110010011	(	adb30110010011,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m100100_0	),
Adb30110010100	(	adb30110010100,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m100100_0	),
Adb30110010101	(	adb30110010101,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m100100_0	),
Adb30110010110	(	adb30110010110,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m100100_0	),
Adb30110010111	(	adb30110010111,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m100100_0	),
Adb30110011000	(	adb30110011000,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m100100_0	),
Adb30110011001	(	adb30110011001,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m100100_0	),
Adb30110011010	(	adb30110011010,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m100100_0	),
Adb30110011011	(	adb30110011011,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m100100_0	),
Adb30110011100	(	adb30110011100,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m100100_0	),
Adb30110011101	(	adb30110011101,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m100100_0	),
Adb30110011110	(	adb30110011110,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m100100_0	),
Adb30110011111	(	adb30110011111,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m100100_0	),
Adb30110100000	(	adb30110100000,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m100100_0	),
Adb30110100001	(	adb30110100001,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m100100_0	),
Adb30110100010	(	adb30110100010,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m100100_0	),
Adb30110100011	(	adb30110100011,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m100100_0	),
Adb30110100100	(	adb30110100100,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m100100_0	),
Adb30110100101	(	adb30110100101,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m100100_0	),
Adb30110100110	(	adb30110100110,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m100100_0	),
Adb30110100111	(	adb30110100111,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m100100_0	),
Adb30110101000	(	adb30110101000,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m100100_0	),
Adb30110101001	(	adb30110101001,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m100100_0	),
Adb30110101010	(	adb30110101010,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m100100_0	),
Adb30110101011	(	adb30110101011,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m100100_0	),
Adb30110101100	(	adb30110101100,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m100100_0	),
Adb30110101101	(	adb30110101101,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m100100_0	),
Adb30110101110	(	adb30110101110,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m100100_0	),
Adb30110101111	(	adb30110101111,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m100100_0	),
Adb30110110000	(	adb30110110000,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m100100_0	),
Adb30110110001	(	adb30110110001,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m100100_0	),
Adb30110110010	(	adb30110110010,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m100100_0	),
Adb30110110011	(	adb30110110011,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m100100_0	),
Adb30110110100	(	adb30110110100,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m100100_0	),
Adb30110110101	(	adb30110110101,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m100100_0	),
Adb30110110110	(	adb30110110110,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m100100_0	),
Adb30110110111	(	adb30110110111,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m100100_0	),
Adb30110111000	(	adb30110111000,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m100100_0	),
Adb30110111001	(	adb30110111001,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m100100_0	),
Adb30110111010	(	adb30110111010,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m100100_0	),
Adb30110111011	(	adb30110111011,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m100100_0	),
Adb30110111100	(	adb30110111100,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m100100_0	),
Adb30110111101	(	adb30110111101,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m100100_0	),
Adb30110111110	(	adb30110111110,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m100100_0	),
Adb30110111111	(	adb30110111111,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m100100_0	),
Adb30111000000	(	adb30111000000,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m100100_0	),
Adb30111000001	(	adb30111000001,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m100100_0	),
Adb30111000010	(	adb30111000010,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m100100_0	),
Adb30111000011	(	adb30111000011,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m100100_0	),
Adb30111000100	(	adb30111000100,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m100100_0	),
Adb30111000101	(	adb30111000101,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m100100_0	),
Adb30111000110	(	adb30111000110,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m100100_0	),
Adb30111000111	(	adb30111000111,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m100100_0	),
Adb30111001000	(	adb30111001000,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m100100_0	),
Adb30111001001	(	adb30111001001,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m100100_0	),
Adb30111001010	(	adb30111001010,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m100100_0	),
Adb30111001011	(	adb30111001011,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m100100_0	),
Adb30111001100	(	adb30111001100,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m100100_0	),
Adb30111001101	(	adb30111001101,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m100100_0	),
Adb30111001110	(	adb30111001110,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m100100_0	),
Adb30111001111	(	adb30111001111,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m100100_0	),
Adb30111010000	(	adb30111010000,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m100100_0	),
Adb30111010001	(	adb30111010001,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m100100_0	),
Adb30111010010	(	adb30111010010,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m100100_0	),
Adb30111010011	(	adb30111010011,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m100100_0	),
Adb30111010100	(	adb30111010100,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m100100_0	),
Adb30111010101	(	adb30111010101,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m100100_0	),
Adb30111010110	(	adb30111010110,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m100100_0	),
Adb30111010111	(	adb30111010111,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m100100_0	),
Adb30111011000	(	adb30111011000,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m100100_0	),
Adb30111011001	(	adb30111011001,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m100100_0	),
Adb30111011010	(	adb30111011010,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m100100_0	),
Adb30111011011	(	adb30111011011,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m100100_0	),
Adb30111011100	(	adb30111011100,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m100100_0	),
Adb30111011101	(	adb30111011101,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m100100_0	),
Adb30111011110	(	adb30111011110,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m100100_0	),
Adb30111011111	(	adb30111011111,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m100100_0	),
Adb30111100000	(	adb30111100000,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m100100_0	),
Adb30111100001	(	adb30111100001,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m100100_0	),
Adb30111100010	(	adb30111100010,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m100100_0	),
Adb30111100011	(	adb30111100011,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m100100_0	),
Adb30111100100	(	adb30111100100,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m100100_0	),
Adb30111100101	(	adb30111100101,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m100100_0	),
Adb30111100110	(	adb30111100110,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m100100_0	),
Adb30111100111	(	adb30111100111,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m100100_0	),
Adb30111101000	(	adb30111101000,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m100100_0	),
Adb30111101001	(	adb30111101001,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m100100_0	),
Adb30111101010	(	adb30111101010,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m100100_0	),
Adb30111101011	(	adb30111101011,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m100100_0	),
Adb30111101100	(	adb30111101100,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m100100_0	),
Adb30111101101	(	adb30111101101,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m100100_0	),
Adb30111101110	(	adb30111101110,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m100100_0	),
Adb30111101111	(	adb30111101111,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m100100_0	),
Adb30111110000	(	adb30111110000,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m100100_0	),
Adb30111110001	(	adb30111110001,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m100100_0	),
Adb30111110010	(	adb30111110010,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m100100_0	),
Adb30111110011	(	adb30111110011,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m100100_0	),
Adb30111110100	(	adb30111110100,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m100100_0	),
Adb30111110101	(	adb30111110101,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m100100_0	),
Adb30111110110	(	adb30111110110,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m100100_0	),
Adb30111110111	(	adb30111110111,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m100100_0	),
Adb30111111000	(	adb30111111000,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m100100_0	),
Adb30111111001	(	adb30111111001,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m100100_0	),
Adb30111111010	(	adb30111111010,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m100100_0	),
Adb30111111011	(	adb30111111011,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m100100_0	),
Adb30111111100	(	adb30111111100,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m100100_0	),
Adb30111111101	(	adb30111111101,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m100100_0	),
Adb30111111110	(	adb30111111110,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m100100_0	),
Adb30111111111	(	adb30111111111,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m100100_0	),
Adb31000000000	(	adb31000000000,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m011100_0	),
Adb31000000001	(	adb31000000001,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m011100_0	),
Adb31000000010	(	adb31000000010,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m011100_0	),
Adb31000000011	(	adb31000000011,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m011100_0	),
Adb31000000100	(	adb31000000100,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m011100_0	),
Adb31000000101	(	adb31000000101,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m011100_0	),
Adb31000000110	(	adb31000000110,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m011100_0	),
Adb31000000111	(	adb31000000111,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m011100_0	),
Adb31000001000	(	adb31000001000,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m011100_0	),
Adb31000001001	(	adb31000001001,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m011100_0	),
Adb31000001010	(	adb31000001010,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m011100_0	),
Adb31000001011	(	adb31000001011,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m011100_0	),
Adb31000001100	(	adb31000001100,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m011100_0	),
Adb31000001101	(	adb31000001101,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m011100_0	),
Adb31000001110	(	adb31000001110,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m011100_0	),
Adb31000001111	(	adb31000001111,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m011100_0	),
Adb31000010000	(	adb31000010000,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m011100_0	),
Adb31000010001	(	adb31000010001,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m011100_0	),
Adb31000010010	(	adb31000010010,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m011100_0	),
Adb31000010011	(	adb31000010011,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m011100_0	),
Adb31000010100	(	adb31000010100,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m011100_0	),
Adb31000010101	(	adb31000010101,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m011100_0	),
Adb31000010110	(	adb31000010110,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m011100_0	),
Adb31000010111	(	adb31000010111,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m011100_0	),
Adb31000011000	(	adb31000011000,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m011100_0	),
Adb31000011001	(	adb31000011001,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m011100_0	),
Adb31000011010	(	adb31000011010,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m011100_0	),
Adb31000011011	(	adb31000011011,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m011100_0	),
Adb31000011100	(	adb31000011100,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m011100_0	),
Adb31000011101	(	adb31000011101,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m011100_0	),
Adb31000011110	(	adb31000011110,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m011100_0	),
Adb31000011111	(	adb31000011111,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m011100_0	),
Adb31000100000	(	adb31000100000,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m011100_0	),
Adb31000100001	(	adb31000100001,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m011100_0	),
Adb31000100010	(	adb31000100010,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m011100_0	),
Adb31000100011	(	adb31000100011,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m011100_0	),
Adb31000100100	(	adb31000100100,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m011100_0	),
Adb31000100101	(	adb31000100101,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m011100_0	),
Adb31000100110	(	adb31000100110,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m011100_0	),
Adb31000100111	(	adb31000100111,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m011100_0	),
Adb31000101000	(	adb31000101000,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m011100_0	),
Adb31000101001	(	adb31000101001,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m011100_0	),
Adb31000101010	(	adb31000101010,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m011100_0	),
Adb31000101011	(	adb31000101011,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m011100_0	),
Adb31000101100	(	adb31000101100,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m011100_0	),
Adb31000101101	(	adb31000101101,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m011100_0	),
Adb31000101110	(	adb31000101110,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m011100_0	),
Adb31000101111	(	adb31000101111,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m011100_0	),
Adb31000110000	(	adb31000110000,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m011100_0	),
Adb31000110001	(	adb31000110001,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m011100_0	),
Adb31000110010	(	adb31000110010,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m011100_0	),
Adb31000110011	(	adb31000110011,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m011100_0	),
Adb31000110100	(	adb31000110100,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m011100_0	),
Adb31000110101	(	adb31000110101,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m011100_0	),
Adb31000110110	(	adb31000110110,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m011100_0	),
Adb31000110111	(	adb31000110111,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m011100_0	),
Adb31000111000	(	adb31000111000,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m011100_0	),
Adb31000111001	(	adb31000111001,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m011100_0	),
Adb31000111010	(	adb31000111010,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m011100_0	),
Adb31000111011	(	adb31000111011,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m011100_0	),
Adb31000111100	(	adb31000111100,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m011100_0	),
Adb31000111101	(	adb31000111101,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m011100_0	),
Adb31000111110	(	adb31000111110,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m011100_0	),
Adb31000111111	(	adb31000111111,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m011100_0	),
Adb31001000000	(	adb31001000000,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m011100_0	),
Adb31001000001	(	adb31001000001,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m011100_0	),
Adb31001000010	(	adb31001000010,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m011100_0	),
Adb31001000011	(	adb31001000011,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m011100_0	),
Adb31001000100	(	adb31001000100,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m011100_0	),
Adb31001000101	(	adb31001000101,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m011100_0	),
Adb31001000110	(	adb31001000110,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m011100_0	),
Adb31001000111	(	adb31001000111,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m011100_0	),
Adb31001001000	(	adb31001001000,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m011100_0	),
Adb31001001001	(	adb31001001001,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m011100_0	),
Adb31001001010	(	adb31001001010,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m011100_0	),
Adb31001001011	(	adb31001001011,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m011100_0	),
Adb31001001100	(	adb31001001100,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m011100_0	),
Adb31001001101	(	adb31001001101,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m011100_0	),
Adb31001001110	(	adb31001001110,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m011100_0	),
Adb31001001111	(	adb31001001111,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m011100_0	),
Adb31001010000	(	adb31001010000,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m011100_0	),
Adb31001010001	(	adb31001010001,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m011100_0	),
Adb31001010010	(	adb31001010010,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m011100_0	),
Adb31001010011	(	adb31001010011,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m011100_0	),
Adb31001010100	(	adb31001010100,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m011100_0	),
Adb31001010101	(	adb31001010101,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m011100_0	),
Adb31001010110	(	adb31001010110,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m011100_0	),
Adb31001010111	(	adb31001010111,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m011100_0	),
Adb31001011000	(	adb31001011000,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m011100_0	),
Adb31001011001	(	adb31001011001,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m011100_0	),
Adb31001011010	(	adb31001011010,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m011100_0	),
Adb31001011011	(	adb31001011011,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m011100_0	),
Adb31001011100	(	adb31001011100,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m011100_0	),
Adb31001011101	(	adb31001011101,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m011100_0	),
Adb31001011110	(	adb31001011110,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m011100_0	),
Adb31001011111	(	adb31001011111,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m011100_0	),
Adb31001100000	(	adb31001100000,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m011100_0	),
Adb31001100001	(	adb31001100001,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m011100_0	),
Adb31001100010	(	adb31001100010,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m011100_0	),
Adb31001100011	(	adb31001100011,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m011100_0	),
Adb31001100100	(	adb31001100100,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m011100_0	),
Adb31001100101	(	adb31001100101,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m011100_0	),
Adb31001100110	(	adb31001100110,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m011100_0	),
Adb31001100111	(	adb31001100111,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m011100_0	),
Adb31001101000	(	adb31001101000,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m011100_0	),
Adb31001101001	(	adb31001101001,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m011100_0	),
Adb31001101010	(	adb31001101010,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m011100_0	),
Adb31001101011	(	adb31001101011,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m011100_0	),
Adb31001101100	(	adb31001101100,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m011100_0	),
Adb31001101101	(	adb31001101101,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m011100_0	),
Adb31001101110	(	adb31001101110,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m011100_0	),
Adb31001101111	(	adb31001101111,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m011100_0	),
Adb31001110000	(	adb31001110000,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m011100_0	),
Adb31001110001	(	adb31001110001,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m011100_0	),
Adb31001110010	(	adb31001110010,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m011100_0	),
Adb31001110011	(	adb31001110011,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m011100_0	),
Adb31001110100	(	adb31001110100,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m011100_0	),
Adb31001110101	(	adb31001110101,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m011100_0	),
Adb31001110110	(	adb31001110110,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m011100_0	),
Adb31001110111	(	adb31001110111,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m011100_0	),
Adb31001111000	(	adb31001111000,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m011100_0	),
Adb31001111001	(	adb31001111001,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m011100_0	),
Adb31001111010	(	adb31001111010,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m011100_0	),
Adb31001111011	(	adb31001111011,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m011100_0	),
Adb31001111100	(	adb31001111100,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m011100_0	),
Adb31001111101	(	adb31001111101,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m011100_0	),
Adb31001111110	(	adb31001111110,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m011100_0	),
Adb31001111111	(	adb31001111111,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m011100_0	),
Adb31010000000	(	adb31010000000,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m010100_0	),
Adb31010000001	(	adb31010000001,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m010100_0	),
Adb31010000010	(	adb31010000010,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m010100_0	),
Adb31010000011	(	adb31010000011,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m010100_0	),
Adb31010000100	(	adb31010000100,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m010100_0	),
Adb31010000101	(	adb31010000101,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m010100_0	),
Adb31010000110	(	adb31010000110,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m010100_0	),
Adb31010000111	(	adb31010000111,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m010100_0	),
Adb31010001000	(	adb31010001000,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m010100_0	),
Adb31010001001	(	adb31010001001,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m010100_0	),
Adb31010001010	(	adb31010001010,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m010100_0	),
Adb31010001011	(	adb31010001011,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m010100_0	),
Adb31010001100	(	adb31010001100,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m010100_0	),
Adb31010001101	(	adb31010001101,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m010100_0	),
Adb31010001110	(	adb31010001110,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m010100_0	),
Adb31010001111	(	adb31010001111,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m010100_0	),
Adb31010010000	(	adb31010010000,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m010100_0	),
Adb31010010001	(	adb31010010001,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m010100_0	),
Adb31010010010	(	adb31010010010,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m010100_0	),
Adb31010010011	(	adb31010010011,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m010100_0	),
Adb31010010100	(	adb31010010100,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m010100_0	),
Adb31010010101	(	adb31010010101,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m010100_0	),
Adb31010010110	(	adb31010010110,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m010100_0	),
Adb31010010111	(	adb31010010111,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m010100_0	),
Adb31010011000	(	adb31010011000,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m010100_0	),
Adb31010011001	(	adb31010011001,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m010100_0	),
Adb31010011010	(	adb31010011010,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m010100_0	),
Adb31010011011	(	adb31010011011,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m010100_0	),
Adb31010011100	(	adb31010011100,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m010100_0	),
Adb31010011101	(	adb31010011101,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m010100_0	),
Adb31010011110	(	adb31010011110,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m010100_0	),
Adb31010011111	(	adb31010011111,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m010100_0	),
Adb31010100000	(	adb31010100000,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m010100_0	),
Adb31010100001	(	adb31010100001,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m010100_0	),
Adb31010100010	(	adb31010100010,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m010100_0	),
Adb31010100011	(	adb31010100011,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m010100_0	),
Adb31010100100	(	adb31010100100,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m010100_0	),
Adb31010100101	(	adb31010100101,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m010100_0	),
Adb31010100110	(	adb31010100110,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m010100_0	),
Adb31010100111	(	adb31010100111,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m010100_0	),
Adb31010101000	(	adb31010101000,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m010100_0	),
Adb31010101001	(	adb31010101001,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m010100_0	),
Adb31010101010	(	adb31010101010,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m010100_0	),
Adb31010101011	(	adb31010101011,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m010100_0	),
Adb31010101100	(	adb31010101100,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m010100_0	),
Adb31010101101	(	adb31010101101,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m010100_0	),
Adb31010101110	(	adb31010101110,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m010100_0	),
Adb31010101111	(	adb31010101111,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m010100_0	),
Adb31010110000	(	adb31010110000,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m010100_0	),
Adb31010110001	(	adb31010110001,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m010100_0	),
Adb31010110010	(	adb31010110010,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m010100_0	),
Adb31010110011	(	adb31010110011,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m010100_0	),
Adb31010110100	(	adb31010110100,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m010100_0	),
Adb31010110101	(	adb31010110101,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m010100_0	),
Adb31010110110	(	adb31010110110,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m010100_0	),
Adb31010110111	(	adb31010110111,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m010100_0	),
Adb31010111000	(	adb31010111000,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m010100_0	),
Adb31010111001	(	adb31010111001,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m010100_0	),
Adb31010111010	(	adb31010111010,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m010100_0	),
Adb31010111011	(	adb31010111011,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m010100_0	),
Adb31010111100	(	adb31010111100,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m010100_0	),
Adb31010111101	(	adb31010111101,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m010100_0	),
Adb31010111110	(	adb31010111110,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m010100_0	),
Adb31010111111	(	adb31010111111,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m010100_0	),
Adb31011000000	(	adb31011000000,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m010100_0	),
Adb31011000001	(	adb31011000001,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m010100_0	),
Adb31011000010	(	adb31011000010,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m010100_0	),
Adb31011000011	(	adb31011000011,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m010100_0	),
Adb31011000100	(	adb31011000100,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m010100_0	),
Adb31011000101	(	adb31011000101,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m010100_0	),
Adb31011000110	(	adb31011000110,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m010100_0	),
Adb31011000111	(	adb31011000111,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m010100_0	),
Adb31011001000	(	adb31011001000,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m010100_0	),
Adb31011001001	(	adb31011001001,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m010100_0	),
Adb31011001010	(	adb31011001010,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m010100_0	),
Adb31011001011	(	adb31011001011,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m010100_0	),
Adb31011001100	(	adb31011001100,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m010100_0	),
Adb31011001101	(	adb31011001101,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m010100_0	),
Adb31011001110	(	adb31011001110,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m010100_0	),
Adb31011001111	(	adb31011001111,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m010100_0	),
Adb31011010000	(	adb31011010000,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m010100_0	),
Adb31011010001	(	adb31011010001,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m010100_0	),
Adb31011010010	(	adb31011010010,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m010100_0	),
Adb31011010011	(	adb31011010011,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m010100_0	),
Adb31011010100	(	adb31011010100,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m010100_0	),
Adb31011010101	(	adb31011010101,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m010100_0	),
Adb31011010110	(	adb31011010110,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m010100_0	),
Adb31011010111	(	adb31011010111,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m010100_0	),
Adb31011011000	(	adb31011011000,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m010100_0	),
Adb31011011001	(	adb31011011001,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m010100_0	),
Adb31011011010	(	adb31011011010,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m010100_0	),
Adb31011011011	(	adb31011011011,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m010100_0	),
Adb31011011100	(	adb31011011100,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m010100_0	),
Adb31011011101	(	adb31011011101,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m010100_0	),
Adb31011011110	(	adb31011011110,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m010100_0	),
Adb31011011111	(	adb31011011111,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m010100_0	),
Adb31011100000	(	adb31011100000,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m010100_0	),
Adb31011100001	(	adb31011100001,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m010100_0	),
Adb31011100010	(	adb31011100010,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m010100_0	),
Adb31011100011	(	adb31011100011,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m010100_0	),
Adb31011100100	(	adb31011100100,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m010100_0	),
Adb31011100101	(	adb31011100101,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m010100_0	),
Adb31011100110	(	adb31011100110,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m010100_0	),
Adb31011100111	(	adb31011100111,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m010100_0	),
Adb31011101000	(	adb31011101000,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m010100_0	),
Adb31011101001	(	adb31011101001,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m010100_0	),
Adb31011101010	(	adb31011101010,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m010100_0	),
Adb31011101011	(	adb31011101011,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m010100_0	),
Adb31011101100	(	adb31011101100,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m010100_0	),
Adb31011101101	(	adb31011101101,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m010100_0	),
Adb31011101110	(	adb31011101110,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m010100_0	),
Adb31011101111	(	adb31011101111,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m010100_0	),
Adb31011110000	(	adb31011110000,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m010100_0	),
Adb31011110001	(	adb31011110001,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m010100_0	),
Adb31011110010	(	adb31011110010,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m010100_0	),
Adb31011110011	(	adb31011110011,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m010100_0	),
Adb31011110100	(	adb31011110100,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m010100_0	),
Adb31011110101	(	adb31011110101,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m010100_0	),
Adb31011110110	(	adb31011110110,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m010100_0	),
Adb31011110111	(	adb31011110111,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m010100_0	),
Adb31011111000	(	adb31011111000,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m010100_0	),
Adb31011111001	(	adb31011111001,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m010100_0	),
Adb31011111010	(	adb31011111010,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m010100_0	),
Adb31011111011	(	adb31011111011,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m010100_0	),
Adb31011111100	(	adb31011111100,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m010100_0	),
Adb31011111101	(	adb31011111101,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m010100_0	),
Adb31011111110	(	adb31011111110,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m010100_0	),
Adb31011111111	(	adb31011111111,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m010100_0	),
Adb31100000000	(	adb31100000000,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m001100_0	),
Adb31100000001	(	adb31100000001,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m001100_0	),
Adb31100000010	(	adb31100000010,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m001100_0	),
Adb31100000011	(	adb31100000011,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m001100_0	),
Adb31100000100	(	adb31100000100,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m001100_0	),
Adb31100000101	(	adb31100000101,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m001100_0	),
Adb31100000110	(	adb31100000110,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m001100_0	),
Adb31100000111	(	adb31100000111,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m001100_0	),
Adb31100001000	(	adb31100001000,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m001100_0	),
Adb31100001001	(	adb31100001001,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m001100_0	),
Adb31100001010	(	adb31100001010,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m001100_0	),
Adb31100001011	(	adb31100001011,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m001100_0	),
Adb31100001100	(	adb31100001100,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m001100_0	),
Adb31100001101	(	adb31100001101,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m001100_0	),
Adb31100001110	(	adb31100001110,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m001100_0	),
Adb31100001111	(	adb31100001111,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m001100_0	),
Adb31100010000	(	adb31100010000,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m001100_0	),
Adb31100010001	(	adb31100010001,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m001100_0	),
Adb31100010010	(	adb31100010010,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m001100_0	),
Adb31100010011	(	adb31100010011,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m001100_0	),
Adb31100010100	(	adb31100010100,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m001100_0	),
Adb31100010101	(	adb31100010101,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m001100_0	),
Adb31100010110	(	adb31100010110,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m001100_0	),
Adb31100010111	(	adb31100010111,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m001100_0	),
Adb31100011000	(	adb31100011000,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m001100_0	),
Adb31100011001	(	adb31100011001,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m001100_0	),
Adb31100011010	(	adb31100011010,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m001100_0	),
Adb31100011011	(	adb31100011011,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m001100_0	),
Adb31100011100	(	adb31100011100,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m001100_0	),
Adb31100011101	(	adb31100011101,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m001100_0	),
Adb31100011110	(	adb31100011110,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m001100_0	),
Adb31100011111	(	adb31100011111,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m001100_0	),
Adb31100100000	(	adb31100100000,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m001100_0	),
Adb31100100001	(	adb31100100001,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m001100_0	),
Adb31100100010	(	adb31100100010,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m001100_0	),
Adb31100100011	(	adb31100100011,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m001100_0	),
Adb31100100100	(	adb31100100100,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m001100_0	),
Adb31100100101	(	adb31100100101,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m001100_0	),
Adb31100100110	(	adb31100100110,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m001100_0	),
Adb31100100111	(	adb31100100111,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m001100_0	),
Adb31100101000	(	adb31100101000,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m001100_0	),
Adb31100101001	(	adb31100101001,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m001100_0	),
Adb31100101010	(	adb31100101010,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m001100_0	),
Adb31100101011	(	adb31100101011,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m001100_0	),
Adb31100101100	(	adb31100101100,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m001100_0	),
Adb31100101101	(	adb31100101101,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m001100_0	),
Adb31100101110	(	adb31100101110,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m001100_0	),
Adb31100101111	(	adb31100101111,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m001100_0	),
Adb31100110000	(	adb31100110000,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m001100_0	),
Adb31100110001	(	adb31100110001,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m001100_0	),
Adb31100110010	(	adb31100110010,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m001100_0	),
Adb31100110011	(	adb31100110011,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m001100_0	),
Adb31100110100	(	adb31100110100,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m001100_0	),
Adb31100110101	(	adb31100110101,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m001100_0	),
Adb31100110110	(	adb31100110110,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m001100_0	),
Adb31100110111	(	adb31100110111,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m001100_0	),
Adb31100111000	(	adb31100111000,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m001100_0	),
Adb31100111001	(	adb31100111001,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m001100_0	),
Adb31100111010	(	adb31100111010,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m001100_0	),
Adb31100111011	(	adb31100111011,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m001100_0	),
Adb31100111100	(	adb31100111100,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m001100_0	),
Adb31100111101	(	adb31100111101,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m001100_0	),
Adb31100111110	(	adb31100111110,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m001100_0	),
Adb31100111111	(	adb31100111111,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m001100_0	),
Adb31101000000	(	adb31101000000,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m001100_0	),
Adb31101000001	(	adb31101000001,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m001100_0	),
Adb31101000010	(	adb31101000010,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m001100_0	),
Adb31101000011	(	adb31101000011,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m001100_0	),
Adb31101000100	(	adb31101000100,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m001100_0	),
Adb31101000101	(	adb31101000101,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m001100_0	),
Adb31101000110	(	adb31101000110,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m001100_0	),
Adb31101000111	(	adb31101000111,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m001100_0	),
Adb31101001000	(	adb31101001000,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m001100_0	),
Adb31101001001	(	adb31101001001,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m001100_0	),
Adb31101001010	(	adb31101001010,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m001100_0	),
Adb31101001011	(	adb31101001011,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m001100_0	),
Adb31101001100	(	adb31101001100,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m001100_0	),
Adb31101001101	(	adb31101001101,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m001100_0	),
Adb31101001110	(	adb31101001110,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m001100_0	),
Adb31101001111	(	adb31101001111,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m001100_0	),
Adb31101010000	(	adb31101010000,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m001100_0	),
Adb31101010001	(	adb31101010001,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m001100_0	),
Adb31101010010	(	adb31101010010,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m001100_0	),
Adb31101010011	(	adb31101010011,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m001100_0	),
Adb31101010100	(	adb31101010100,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m001100_0	),
Adb31101010101	(	adb31101010101,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m001100_0	),
Adb31101010110	(	adb31101010110,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m001100_0	),
Adb31101010111	(	adb31101010111,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m001100_0	),
Adb31101011000	(	adb31101011000,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m001100_0	),
Adb31101011001	(	adb31101011001,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m001100_0	),
Adb31101011010	(	adb31101011010,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m001100_0	),
Adb31101011011	(	adb31101011011,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m001100_0	),
Adb31101011100	(	adb31101011100,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m001100_0	),
Adb31101011101	(	adb31101011101,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m001100_0	),
Adb31101011110	(	adb31101011110,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m001100_0	),
Adb31101011111	(	adb31101011111,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m001100_0	),
Adb31101100000	(	adb31101100000,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m001100_0	),
Adb31101100001	(	adb31101100001,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m001100_0	),
Adb31101100010	(	adb31101100010,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m001100_0	),
Adb31101100011	(	adb31101100011,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m001100_0	),
Adb31101100100	(	adb31101100100,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m001100_0	),
Adb31101100101	(	adb31101100101,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m001100_0	),
Adb31101100110	(	adb31101100110,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m001100_0	),
Adb31101100111	(	adb31101100111,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m001100_0	),
Adb31101101000	(	adb31101101000,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m001100_0	),
Adb31101101001	(	adb31101101001,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m001100_0	),
Adb31101101010	(	adb31101101010,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m001100_0	),
Adb31101101011	(	adb31101101011,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m001100_0	),
Adb31101101100	(	adb31101101100,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m001100_0	),
Adb31101101101	(	adb31101101101,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m001100_0	),
Adb31101101110	(	adb31101101110,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m001100_0	),
Adb31101101111	(	adb31101101111,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m001100_0	),
Adb31101110000	(	adb31101110000,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m001100_0	),
Adb31101110001	(	adb31101110001,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m001100_0	),
Adb31101110010	(	adb31101110010,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m001100_0	),
Adb31101110011	(	adb31101110011,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m001100_0	),
Adb31101110100	(	adb31101110100,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m001100_0	),
Adb31101110101	(	adb31101110101,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m001100_0	),
Adb31101110110	(	adb31101110110,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m001100_0	),
Adb31101110111	(	adb31101110111,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m001100_0	),
Adb31101111000	(	adb31101111000,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m001100_0	),
Adb31101111001	(	adb31101111001,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m001100_0	),
Adb31101111010	(	adb31101111010,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m001100_0	),
Adb31101111011	(	adb31101111011,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m001100_0	),
Adb31101111100	(	adb31101111100,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m001100_0	),
Adb31101111101	(	adb31101111101,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m001100_0	),
Adb31101111110	(	adb31101111110,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m001100_0	),
Adb31101111111	(	adb31101111111,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m001100_0	),
Adb31110000000	(	adb31110000000,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m000100_0	),
Adb31110000001	(	adb31110000001,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m000100_0	),
Adb31110000010	(	adb31110000010,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m000100_0	),
Adb31110000011	(	adb31110000011,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m000100_0	),
Adb31110000100	(	adb31110000100,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m000100_0	),
Adb31110000101	(	adb31110000101,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m000100_0	),
Adb31110000110	(	adb31110000110,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m000100_0	),
Adb31110000111	(	adb31110000111,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m000100_0	),
Adb31110001000	(	adb31110001000,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m000100_0	),
Adb31110001001	(	adb31110001001,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m000100_0	),
Adb31110001010	(	adb31110001010,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m000100_0	),
Adb31110001011	(	adb31110001011,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m000100_0	),
Adb31110001100	(	adb31110001100,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m000100_0	),
Adb31110001101	(	adb31110001101,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m000100_0	),
Adb31110001110	(	adb31110001110,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m000100_0	),
Adb31110001111	(	adb31110001111,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m000100_0	),
Adb31110010000	(	adb31110010000,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m000100_0	),
Adb31110010001	(	adb31110010001,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m000100_0	),
Adb31110010010	(	adb31110010010,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m000100_0	),
Adb31110010011	(	adb31110010011,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m000100_0	),
Adb31110010100	(	adb31110010100,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m000100_0	),
Adb31110010101	(	adb31110010101,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m000100_0	),
Adb31110010110	(	adb31110010110,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m000100_0	),
Adb31110010111	(	adb31110010111,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m000100_0	),
Adb31110011000	(	adb31110011000,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m000100_0	),
Adb31110011001	(	adb31110011001,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m000100_0	),
Adb31110011010	(	adb31110011010,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m000100_0	),
Adb31110011011	(	adb31110011011,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m000100_0	),
Adb31110011100	(	adb31110011100,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m000100_0	),
Adb31110011101	(	adb31110011101,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m000100_0	),
Adb31110011110	(	adb31110011110,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m000100_0	),
Adb31110011111	(	adb31110011111,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m000100_0	),
Adb31110100000	(	adb31110100000,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m000100_0	),
Adb31110100001	(	adb31110100001,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m000100_0	),
Adb31110100010	(	adb31110100010,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m000100_0	),
Adb31110100011	(	adb31110100011,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m000100_0	),
Adb31110100100	(	adb31110100100,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m000100_0	),
Adb31110100101	(	adb31110100101,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m000100_0	),
Adb31110100110	(	adb31110100110,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m000100_0	),
Adb31110100111	(	adb31110100111,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m000100_0	),
Adb31110101000	(	adb31110101000,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m000100_0	),
Adb31110101001	(	adb31110101001,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m000100_0	),
Adb31110101010	(	adb31110101010,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m000100_0	),
Adb31110101011	(	adb31110101011,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m000100_0	),
Adb31110101100	(	adb31110101100,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m000100_0	),
Adb31110101101	(	adb31110101101,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m000100_0	),
Adb31110101110	(	adb31110101110,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m000100_0	),
Adb31110101111	(	adb31110101111,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m000100_0	),
Adb31110110000	(	adb31110110000,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m000100_0	),
Adb31110110001	(	adb31110110001,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m000100_0	),
Adb31110110010	(	adb31110110010,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m000100_0	),
Adb31110110011	(	adb31110110011,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m000100_0	),
Adb31110110100	(	adb31110110100,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m000100_0	),
Adb31110110101	(	adb31110110101,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m000100_0	),
Adb31110110110	(	adb31110110110,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m000100_0	),
Adb31110110111	(	adb31110110111,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m000100_0	),
Adb31110111000	(	adb31110111000,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m000100_0	),
Adb31110111001	(	adb31110111001,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m000100_0	),
Adb31110111010	(	adb31110111010,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m000100_0	),
Adb31110111011	(	adb31110111011,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m000100_0	),
Adb31110111100	(	adb31110111100,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m000100_0	),
Adb31110111101	(	adb31110111101,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m000100_0	),
Adb31110111110	(	adb31110111110,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m000100_0	),
Adb31110111111	(	adb31110111111,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m000100_0	),
Adb31111000000	(	adb31111000000,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m000100_0	),
Adb31111000001	(	adb31111000001,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m000100_0	),
Adb31111000010	(	adb31111000010,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m000100_0	),
Adb31111000011	(	adb31111000011,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m000100_0	),
Adb31111000100	(	adb31111000100,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m000100_0	),
Adb31111000101	(	adb31111000101,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m000100_0	),
Adb31111000110	(	adb31111000110,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m000100_0	),
Adb31111000111	(	adb31111000111,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m000100_0	),
Adb31111001000	(	adb31111001000,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m000100_0	),
Adb31111001001	(	adb31111001001,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m000100_0	),
Adb31111001010	(	adb31111001010,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m000100_0	),
Adb31111001011	(	adb31111001011,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m000100_0	),
Adb31111001100	(	adb31111001100,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m000100_0	),
Adb31111001101	(	adb31111001101,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m000100_0	),
Adb31111001110	(	adb31111001110,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m000100_0	),
Adb31111001111	(	adb31111001111,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m000100_0	),
Adb31111010000	(	adb31111010000,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m000100_0	),
Adb31111010001	(	adb31111010001,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m000100_0	),
Adb31111010010	(	adb31111010010,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m000100_0	),
Adb31111010011	(	adb31111010011,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m000100_0	),
Adb31111010100	(	adb31111010100,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m000100_0	),
Adb31111010101	(	adb31111010101,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m000100_0	),
Adb31111010110	(	adb31111010110,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m000100_0	),
Adb31111010111	(	adb31111010111,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m000100_0	),
Adb31111011000	(	adb31111011000,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m000100_0	),
Adb31111011001	(	adb31111011001,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m000100_0	),
Adb31111011010	(	adb31111011010,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m000100_0	),
Adb31111011011	(	adb31111011011,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m000100_0	),
Adb31111011100	(	adb31111011100,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m000100_0	),
Adb31111011101	(	adb31111011101,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m000100_0	),
Adb31111011110	(	adb31111011110,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m000100_0	),
Adb31111011111	(	adb31111011111,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m000100_0	),
Adb31111100000	(	adb31111100000,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m000100_0	),
Adb31111100001	(	adb31111100001,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m000100_0	),
Adb31111100010	(	adb31111100010,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m000100_0	),
Adb31111100011	(	adb31111100011,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m000100_0	),
Adb31111100100	(	adb31111100100,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m000100_0	),
Adb31111100101	(	adb31111100101,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m000100_0	),
Adb31111100110	(	adb31111100110,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m000100_0	),
Adb31111100111	(	adb31111100111,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m000100_0	),
Adb31111101000	(	adb31111101000,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m000100_0	),
Adb31111101001	(	adb31111101001,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m000100_0	),
Adb31111101010	(	adb31111101010,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m000100_0	),
Adb31111101011	(	adb31111101011,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m000100_0	),
Adb31111101100	(	adb31111101100,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m000100_0	),
Adb31111101101	(	adb31111101101,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m000100_0	),
Adb31111101110	(	adb31111101110,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m000100_0	),
Adb31111101111	(	adb31111101111,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m000100_0	),
Adb31111110000	(	adb31111110000,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m000100_0	),
Adb31111110001	(	adb31111110001,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m000100_0	),
Adb31111110010	(	adb31111110010,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m000100_0	),
Adb31111110011	(	adb31111110011,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m000100_0	),
Adb31111110100	(	adb31111110100,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m000100_0	),
Adb31111110101	(	adb31111110101,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m000100_0	),
Adb31111110110	(	adb31111110110,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m000100_0	),
Adb31111110111	(	adb31111110111,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m000100_0	),
Adb31111111000	(	adb31111111000,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m000100_0	),
Adb31111111001	(	adb31111111001,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m000100_0	),
Adb31111111010	(	adb31111111010,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m000100_0	),
Adb31111111011	(	adb31111111011,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m000100_0	),
Adb31111111100	(	adb31111111100,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m000100_0	),
Adb31111111101	(	adb31111111101,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m000100_0	),
Adb31111111110	(	adb31111111110,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m000100_0	),
Adb31111111111	(	adb31111111111,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m000100_0	),
       Adb400(adb400,n0011,n0010,n0009,dbv1),
       Adb401(adb401,n0011,n0010,m0009,m0014),
       Adb410(adb410,n0011,m0010,n0009,dbv1),
       Adb411(adb411,n0011,m0010,m0009,dbv0),
Adb40000000000	(	adb40000000000,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m111011_0	),
Adb40000000001	(	adb40000000001,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m111011_0	),
Adb40000000010	(	adb40000000010,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m111011_0	),
Adb40000000011	(	adb40000000011,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m111011_0	),
Adb40000000100	(	adb40000000100,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m111011_0	),
Adb40000000101	(	adb40000000101,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m111011_0	),
Adb40000000110	(	adb40000000110,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m111011_0	),
Adb40000000111	(	adb40000000111,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m111011_0	),
Adb40000001000	(	adb40000001000,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m111011_0	),
Adb40000001001	(	adb40000001001,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m111011_0	),
Adb40000001010	(	adb40000001010,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m111011_0	),
Adb40000001011	(	adb40000001011,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m111011_0	),
Adb40000001100	(	adb40000001100,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m111011_0	),
Adb40000001101	(	adb40000001101,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m111011_0	),
Adb40000001110	(	adb40000001110,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m111011_0	),
Adb40000001111	(	adb40000001111,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m111011_0	),
Adb40000010000	(	adb40000010000,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m111011_0	),
Adb40000010001	(	adb40000010001,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m111011_0	),
Adb40000010010	(	adb40000010010,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m111011_0	),
Adb40000010011	(	adb40000010011,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m111011_0	),
Adb40000010100	(	adb40000010100,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m111011_0	),
Adb40000010101	(	adb40000010101,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m111011_0	),
Adb40000010110	(	adb40000010110,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m111011_0	),
Adb40000010111	(	adb40000010111,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m111011_0	),
Adb40000011000	(	adb40000011000,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m111011_0	),
Adb40000011001	(	adb40000011001,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m111011_0	),
Adb40000011010	(	adb40000011010,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m111011_0	),
Adb40000011011	(	adb40000011011,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m111011_0	),
Adb40000011100	(	adb40000011100,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m111011_0	),
Adb40000011101	(	adb40000011101,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m111011_0	),
Adb40000011110	(	adb40000011110,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m111011_0	),
Adb40000011111	(	adb40000011111,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m111011_0	),
Adb40000100000	(	adb40000100000,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m111011_0	),
Adb40000100001	(	adb40000100001,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m111011_0	),
Adb40000100010	(	adb40000100010,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m111011_0	),
Adb40000100011	(	adb40000100011,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m111011_0	),
Adb40000100100	(	adb40000100100,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m111011_0	),
Adb40000100101	(	adb40000100101,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m111011_0	),
Adb40000100110	(	adb40000100110,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m111011_0	),
Adb40000100111	(	adb40000100111,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m111011_0	),
Adb40000101000	(	adb40000101000,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m111011_0	),
Adb40000101001	(	adb40000101001,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m111011_0	),
Adb40000101010	(	adb40000101010,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m111011_0	),
Adb40000101011	(	adb40000101011,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m111011_0	),
Adb40000101100	(	adb40000101100,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m111011_0	),
Adb40000101101	(	adb40000101101,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m111011_0	),
Adb40000101110	(	adb40000101110,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m111011_0	),
Adb40000101111	(	adb40000101111,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m111011_0	),
Adb40000110000	(	adb40000110000,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m111011_0	),
Adb40000110001	(	adb40000110001,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m111011_0	),
Adb40000110010	(	adb40000110010,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m111011_0	),
Adb40000110011	(	adb40000110011,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m111011_0	),
Adb40000110100	(	adb40000110100,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m111011_0	),
Adb40000110101	(	adb40000110101,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m111011_0	),
Adb40000110110	(	adb40000110110,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m111011_0	),
Adb40000110111	(	adb40000110111,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m111011_0	),
Adb40000111000	(	adb40000111000,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m111011_0	),
Adb40000111001	(	adb40000111001,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m111011_0	),
Adb40000111010	(	adb40000111010,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m111011_0	),
Adb40000111011	(	adb40000111011,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m111011_0	),
Adb40000111100	(	adb40000111100,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m111011_0	),
Adb40000111101	(	adb40000111101,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m111011_0	),
Adb40000111110	(	adb40000111110,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m111011_0	),
Adb40000111111	(	adb40000111111,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m111011_0	),
Adb40001000000	(	adb40001000000,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m111011_0	),
Adb40001000001	(	adb40001000001,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m111011_0	),
Adb40001000010	(	adb40001000010,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m111011_0	),
Adb40001000011	(	adb40001000011,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m111011_0	),
Adb40001000100	(	adb40001000100,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m111011_0	),
Adb40001000101	(	adb40001000101,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m111011_0	),
Adb40001000110	(	adb40001000110,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m111011_0	),
Adb40001000111	(	adb40001000111,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m111011_0	),
Adb40001001000	(	adb40001001000,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m111011_0	),
Adb40001001001	(	adb40001001001,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m111011_0	),
Adb40001001010	(	adb40001001010,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m111011_0	),
Adb40001001011	(	adb40001001011,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m111011_0	),
Adb40001001100	(	adb40001001100,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m111011_0	),
Adb40001001101	(	adb40001001101,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m111011_0	),
Adb40001001110	(	adb40001001110,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m111011_0	),
Adb40001001111	(	adb40001001111,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m111011_0	),
Adb40001010000	(	adb40001010000,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m111011_0	),
Adb40001010001	(	adb40001010001,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m111011_0	),
Adb40001010010	(	adb40001010010,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m111011_0	),
Adb40001010011	(	adb40001010011,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m111011_0	),
Adb40001010100	(	adb40001010100,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m111011_0	),
Adb40001010101	(	adb40001010101,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m111011_0	),
Adb40001010110	(	adb40001010110,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m111011_0	),
Adb40001010111	(	adb40001010111,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m111011_0	),
Adb40001011000	(	adb40001011000,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m111011_0	),
Adb40001011001	(	adb40001011001,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m111011_0	),
Adb40001011010	(	adb40001011010,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m111011_0	),
Adb40001011011	(	adb40001011011,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m111011_0	),
Adb40001011100	(	adb40001011100,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m111011_0	),
Adb40001011101	(	adb40001011101,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m111011_0	),
Adb40001011110	(	adb40001011110,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m111011_0	),
Adb40001011111	(	adb40001011111,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m111011_0	),
Adb40001100000	(	adb40001100000,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m111011_0	),
Adb40001100001	(	adb40001100001,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m111011_0	),
Adb40001100010	(	adb40001100010,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m111011_0	),
Adb40001100011	(	adb40001100011,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m111011_0	),
Adb40001100100	(	adb40001100100,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m111011_0	),
Adb40001100101	(	adb40001100101,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m111011_0	),
Adb40001100110	(	adb40001100110,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m111011_0	),
Adb40001100111	(	adb40001100111,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m111011_0	),
Adb40001101000	(	adb40001101000,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m111011_0	),
Adb40001101001	(	adb40001101001,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m111011_0	),
Adb40001101010	(	adb40001101010,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m111011_0	),
Adb40001101011	(	adb40001101011,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m111011_0	),
Adb40001101100	(	adb40001101100,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m111011_0	),
Adb40001101101	(	adb40001101101,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m111011_0	),
Adb40001101110	(	adb40001101110,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m111011_0	),
Adb40001101111	(	adb40001101111,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m111011_0	),
Adb40001110000	(	adb40001110000,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m111011_0	),
Adb40001110001	(	adb40001110001,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m111011_0	),
Adb40001110010	(	adb40001110010,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m111011_0	),
Adb40001110011	(	adb40001110011,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m111011_0	),
Adb40001110100	(	adb40001110100,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m111011_0	),
Adb40001110101	(	adb40001110101,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m111011_0	),
Adb40001110110	(	adb40001110110,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m111011_0	),
Adb40001110111	(	adb40001110111,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m111011_0	),
Adb40001111000	(	adb40001111000,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m111011_0	),
Adb40001111001	(	adb40001111001,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m111011_0	),
Adb40001111010	(	adb40001111010,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m111011_0	),
Adb40001111011	(	adb40001111011,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m111011_0	),
Adb40001111100	(	adb40001111100,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m111011_0	),
Adb40001111101	(	adb40001111101,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m111011_0	),
Adb40001111110	(	adb40001111110,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m111011_0	),
Adb40001111111	(	adb40001111111,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m111011_0	),
Adb40010000000	(	adb40010000000,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m110011_0	),
Adb40010000001	(	adb40010000001,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m110011_0	),
Adb40010000010	(	adb40010000010,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m110011_0	),
Adb40010000011	(	adb40010000011,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m110011_0	),
Adb40010000100	(	adb40010000100,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m110011_0	),
Adb40010000101	(	adb40010000101,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m110011_0	),
Adb40010000110	(	adb40010000110,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m110011_0	),
Adb40010000111	(	adb40010000111,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m110011_0	),
Adb40010001000	(	adb40010001000,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m110011_0	),
Adb40010001001	(	adb40010001001,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m110011_0	),
Adb40010001010	(	adb40010001010,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m110011_0	),
Adb40010001011	(	adb40010001011,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m110011_0	),
Adb40010001100	(	adb40010001100,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m110011_0	),
Adb40010001101	(	adb40010001101,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m110011_0	),
Adb40010001110	(	adb40010001110,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m110011_0	),
Adb40010001111	(	adb40010001111,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m110011_0	),
Adb40010010000	(	adb40010010000,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m110011_0	),
Adb40010010001	(	adb40010010001,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m110011_0	),
Adb40010010010	(	adb40010010010,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m110011_0	),
Adb40010010011	(	adb40010010011,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m110011_0	),
Adb40010010100	(	adb40010010100,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m110011_0	),
Adb40010010101	(	adb40010010101,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m110011_0	),
Adb40010010110	(	adb40010010110,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m110011_0	),
Adb40010010111	(	adb40010010111,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m110011_0	),
Adb40010011000	(	adb40010011000,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m110011_0	),
Adb40010011001	(	adb40010011001,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m110011_0	),
Adb40010011010	(	adb40010011010,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m110011_0	),
Adb40010011011	(	adb40010011011,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m110011_0	),
Adb40010011100	(	adb40010011100,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m110011_0	),
Adb40010011101	(	adb40010011101,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m110011_0	),
Adb40010011110	(	adb40010011110,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m110011_0	),
Adb40010011111	(	adb40010011111,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m110011_0	),
Adb40010100000	(	adb40010100000,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m110011_0	),
Adb40010100001	(	adb40010100001,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m110011_0	),
Adb40010100010	(	adb40010100010,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m110011_0	),
Adb40010100011	(	adb40010100011,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m110011_0	),
Adb40010100100	(	adb40010100100,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m110011_0	),
Adb40010100101	(	adb40010100101,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m110011_0	),
Adb40010100110	(	adb40010100110,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m110011_0	),
Adb40010100111	(	adb40010100111,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m110011_0	),
Adb40010101000	(	adb40010101000,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m110011_0	),
Adb40010101001	(	adb40010101001,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m110011_0	),
Adb40010101010	(	adb40010101010,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m110011_0	),
Adb40010101011	(	adb40010101011,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m110011_0	),
Adb40010101100	(	adb40010101100,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m110011_0	),
Adb40010101101	(	adb40010101101,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m110011_0	),
Adb40010101110	(	adb40010101110,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m110011_0	),
Adb40010101111	(	adb40010101111,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m110011_0	),
Adb40010110000	(	adb40010110000,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m110011_0	),
Adb40010110001	(	adb40010110001,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m110011_0	),
Adb40010110010	(	adb40010110010,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m110011_0	),
Adb40010110011	(	adb40010110011,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m110011_0	),
Adb40010110100	(	adb40010110100,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m110011_0	),
Adb40010110101	(	adb40010110101,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m110011_0	),
Adb40010110110	(	adb40010110110,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m110011_0	),
Adb40010110111	(	adb40010110111,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m110011_0	),
Adb40010111000	(	adb40010111000,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m110011_0	),
Adb40010111001	(	adb40010111001,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m110011_0	),
Adb40010111010	(	adb40010111010,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m110011_0	),
Adb40010111011	(	adb40010111011,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m110011_0	),
Adb40010111100	(	adb40010111100,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m110011_0	),
Adb40010111101	(	adb40010111101,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m110011_0	),
Adb40010111110	(	adb40010111110,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m110011_0	),
Adb40010111111	(	adb40010111111,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m110011_0	),
Adb40011000000	(	adb40011000000,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m110011_0	),
Adb40011000001	(	adb40011000001,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m110011_0	),
Adb40011000010	(	adb40011000010,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m110011_0	),
Adb40011000011	(	adb40011000011,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m110011_0	),
Adb40011000100	(	adb40011000100,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m110011_0	),
Adb40011000101	(	adb40011000101,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m110011_0	),
Adb40011000110	(	adb40011000110,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m110011_0	),
Adb40011000111	(	adb40011000111,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m110011_0	),
Adb40011001000	(	adb40011001000,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m110011_0	),
Adb40011001001	(	adb40011001001,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m110011_0	),
Adb40011001010	(	adb40011001010,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m110011_0	),
Adb40011001011	(	adb40011001011,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m110011_0	),
Adb40011001100	(	adb40011001100,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m110011_0	),
Adb40011001101	(	adb40011001101,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m110011_0	),
Adb40011001110	(	adb40011001110,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m110011_0	),
Adb40011001111	(	adb40011001111,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m110011_0	),
Adb40011010000	(	adb40011010000,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m110011_0	),
Adb40011010001	(	adb40011010001,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m110011_0	),
Adb40011010010	(	adb40011010010,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m110011_0	),
Adb40011010011	(	adb40011010011,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m110011_0	),
Adb40011010100	(	adb40011010100,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m110011_0	),
Adb40011010101	(	adb40011010101,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m110011_0	),
Adb40011010110	(	adb40011010110,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m110011_0	),
Adb40011010111	(	adb40011010111,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m110011_0	),
Adb40011011000	(	adb40011011000,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m110011_0	),
Adb40011011001	(	adb40011011001,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m110011_0	),
Adb40011011010	(	adb40011011010,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m110011_0	),
Adb40011011011	(	adb40011011011,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m110011_0	),
Adb40011011100	(	adb40011011100,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m110011_0	),
Adb40011011101	(	adb40011011101,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m110011_0	),
Adb40011011110	(	adb40011011110,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m110011_0	),
Adb40011011111	(	adb40011011111,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m110011_0	),
Adb40011100000	(	adb40011100000,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m110011_0	),
Adb40011100001	(	adb40011100001,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m110011_0	),
Adb40011100010	(	adb40011100010,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m110011_0	),
Adb40011100011	(	adb40011100011,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m110011_0	),
Adb40011100100	(	adb40011100100,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m110011_0	),
Adb40011100101	(	adb40011100101,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m110011_0	),
Adb40011100110	(	adb40011100110,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m110011_0	),
Adb40011100111	(	adb40011100111,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m110011_0	),
Adb40011101000	(	adb40011101000,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m110011_0	),
Adb40011101001	(	adb40011101001,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m110011_0	),
Adb40011101010	(	adb40011101010,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m110011_0	),
Adb40011101011	(	adb40011101011,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m110011_0	),
Adb40011101100	(	adb40011101100,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m110011_0	),
Adb40011101101	(	adb40011101101,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m110011_0	),
Adb40011101110	(	adb40011101110,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m110011_0	),
Adb40011101111	(	adb40011101111,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m110011_0	),
Adb40011110000	(	adb40011110000,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m110011_0	),
Adb40011110001	(	adb40011110001,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m110011_0	),
Adb40011110010	(	adb40011110010,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m110011_0	),
Adb40011110011	(	adb40011110011,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m110011_0	),
Adb40011110100	(	adb40011110100,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m110011_0	),
Adb40011110101	(	adb40011110101,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m110011_0	),
Adb40011110110	(	adb40011110110,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m110011_0	),
Adb40011110111	(	adb40011110111,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m110011_0	),
Adb40011111000	(	adb40011111000,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m110011_0	),
Adb40011111001	(	adb40011111001,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m110011_0	),
Adb40011111010	(	adb40011111010,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m110011_0	),
Adb40011111011	(	adb40011111011,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m110011_0	),
Adb40011111100	(	adb40011111100,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m110011_0	),
Adb40011111101	(	adb40011111101,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m110011_0	),
Adb40011111110	(	adb40011111110,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m110011_0	),
Adb40011111111	(	adb40011111111,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m110011_0	),
Adb40100000000	(	adb40100000000,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m101011_0	),
Adb40100000001	(	adb40100000001,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m101011_0	),
Adb40100000010	(	adb40100000010,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m101011_0	),
Adb40100000011	(	adb40100000011,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m101011_0	),
Adb40100000100	(	adb40100000100,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m101011_0	),
Adb40100000101	(	adb40100000101,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m101011_0	),
Adb40100000110	(	adb40100000110,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m101011_0	),
Adb40100000111	(	adb40100000111,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m101011_0	),
Adb40100001000	(	adb40100001000,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m101011_0	),
Adb40100001001	(	adb40100001001,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m101011_0	),
Adb40100001010	(	adb40100001010,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m101011_0	),
Adb40100001011	(	adb40100001011,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m101011_0	),
Adb40100001100	(	adb40100001100,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m101011_0	),
Adb40100001101	(	adb40100001101,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m101011_0	),
Adb40100001110	(	adb40100001110,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m101011_0	),
Adb40100001111	(	adb40100001111,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m101011_0	),
Adb40100010000	(	adb40100010000,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m101011_0	),
Adb40100010001	(	adb40100010001,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m101011_0	),
Adb40100010010	(	adb40100010010,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m101011_0	),
Adb40100010011	(	adb40100010011,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m101011_0	),
Adb40100010100	(	adb40100010100,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m101011_0	),
Adb40100010101	(	adb40100010101,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m101011_0	),
Adb40100010110	(	adb40100010110,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m101011_0	),
Adb40100010111	(	adb40100010111,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m101011_0	),
Adb40100011000	(	adb40100011000,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m101011_0	),
Adb40100011001	(	adb40100011001,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m101011_0	),
Adb40100011010	(	adb40100011010,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m101011_0	),
Adb40100011011	(	adb40100011011,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m101011_0	),
Adb40100011100	(	adb40100011100,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m101011_0	),
Adb40100011101	(	adb40100011101,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m101011_0	),
Adb40100011110	(	adb40100011110,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m101011_0	),
Adb40100011111	(	adb40100011111,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m101011_0	),
Adb40100100000	(	adb40100100000,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m101011_0	),
Adb40100100001	(	adb40100100001,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m101011_0	),
Adb40100100010	(	adb40100100010,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m101011_0	),
Adb40100100011	(	adb40100100011,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m101011_0	),
Adb40100100100	(	adb40100100100,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m101011_0	),
Adb40100100101	(	adb40100100101,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m101011_0	),
Adb40100100110	(	adb40100100110,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m101011_0	),
Adb40100100111	(	adb40100100111,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m101011_0	),
Adb40100101000	(	adb40100101000,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m101011_0	),
Adb40100101001	(	adb40100101001,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m101011_0	),
Adb40100101010	(	adb40100101010,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m101011_0	),
Adb40100101011	(	adb40100101011,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m101011_0	),
Adb40100101100	(	adb40100101100,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m101011_0	),
Adb40100101101	(	adb40100101101,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m101011_0	),
Adb40100101110	(	adb40100101110,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m101011_0	),
Adb40100101111	(	adb40100101111,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m101011_0	),
Adb40100110000	(	adb40100110000,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m101011_0	),
Adb40100110001	(	adb40100110001,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m101011_0	),
Adb40100110010	(	adb40100110010,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m101011_0	),
Adb40100110011	(	adb40100110011,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m101011_0	),
Adb40100110100	(	adb40100110100,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m101011_0	),
Adb40100110101	(	adb40100110101,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m101011_0	),
Adb40100110110	(	adb40100110110,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m101011_0	),
Adb40100110111	(	adb40100110111,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m101011_0	),
Adb40100111000	(	adb40100111000,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m101011_0	),
Adb40100111001	(	adb40100111001,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m101011_0	),
Adb40100111010	(	adb40100111010,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m101011_0	),
Adb40100111011	(	adb40100111011,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m101011_0	),
Adb40100111100	(	adb40100111100,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m101011_0	),
Adb40100111101	(	adb40100111101,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m101011_0	),
Adb40100111110	(	adb40100111110,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m101011_0	),
Adb40100111111	(	adb40100111111,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m101011_0	),
Adb40101000000	(	adb40101000000,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m101011_0	),
Adb40101000001	(	adb40101000001,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m101011_0	),
Adb40101000010	(	adb40101000010,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m101011_0	),
Adb40101000011	(	adb40101000011,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m101011_0	),
Adb40101000100	(	adb40101000100,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m101011_0	),
Adb40101000101	(	adb40101000101,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m101011_0	),
Adb40101000110	(	adb40101000110,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m101011_0	),
Adb40101000111	(	adb40101000111,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m101011_0	),
Adb40101001000	(	adb40101001000,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m101011_0	),
Adb40101001001	(	adb40101001001,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m101011_0	),
Adb40101001010	(	adb40101001010,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m101011_0	),
Adb40101001011	(	adb40101001011,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m101011_0	),
Adb40101001100	(	adb40101001100,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m101011_0	),
Adb40101001101	(	adb40101001101,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m101011_0	),
Adb40101001110	(	adb40101001110,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m101011_0	),
Adb40101001111	(	adb40101001111,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m101011_0	),
Adb40101010000	(	adb40101010000,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m101011_0	),
Adb40101010001	(	adb40101010001,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m101011_0	),
Adb40101010010	(	adb40101010010,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m101011_0	),
Adb40101010011	(	adb40101010011,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m101011_0	),
Adb40101010100	(	adb40101010100,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m101011_0	),
Adb40101010101	(	adb40101010101,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m101011_0	),
Adb40101010110	(	adb40101010110,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m101011_0	),
Adb40101010111	(	adb40101010111,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m101011_0	),
Adb40101011000	(	adb40101011000,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m101011_0	),
Adb40101011001	(	adb40101011001,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m101011_0	),
Adb40101011010	(	adb40101011010,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m101011_0	),
Adb40101011011	(	adb40101011011,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m101011_0	),
Adb40101011100	(	adb40101011100,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m101011_0	),
Adb40101011101	(	adb40101011101,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m101011_0	),
Adb40101011110	(	adb40101011110,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m101011_0	),
Adb40101011111	(	adb40101011111,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m101011_0	),
Adb40101100000	(	adb40101100000,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m101011_0	),
Adb40101100001	(	adb40101100001,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m101011_0	),
Adb40101100010	(	adb40101100010,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m101011_0	),
Adb40101100011	(	adb40101100011,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m101011_0	),
Adb40101100100	(	adb40101100100,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m101011_0	),
Adb40101100101	(	adb40101100101,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m101011_0	),
Adb40101100110	(	adb40101100110,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m101011_0	),
Adb40101100111	(	adb40101100111,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m101011_0	),
Adb40101101000	(	adb40101101000,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m101011_0	),
Adb40101101001	(	adb40101101001,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m101011_0	),
Adb40101101010	(	adb40101101010,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m101011_0	),
Adb40101101011	(	adb40101101011,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m101011_0	),
Adb40101101100	(	adb40101101100,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m101011_0	),
Adb40101101101	(	adb40101101101,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m101011_0	),
Adb40101101110	(	adb40101101110,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m101011_0	),
Adb40101101111	(	adb40101101111,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m101011_0	),
Adb40101110000	(	adb40101110000,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m101011_0	),
Adb40101110001	(	adb40101110001,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m101011_0	),
Adb40101110010	(	adb40101110010,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m101011_0	),
Adb40101110011	(	adb40101110011,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m101011_0	),
Adb40101110100	(	adb40101110100,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m101011_0	),
Adb40101110101	(	adb40101110101,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m101011_0	),
Adb40101110110	(	adb40101110110,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m101011_0	),
Adb40101110111	(	adb40101110111,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m101011_0	),
Adb40101111000	(	adb40101111000,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m101011_0	),
Adb40101111001	(	adb40101111001,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m101011_0	),
Adb40101111010	(	adb40101111010,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m101011_0	),
Adb40101111011	(	adb40101111011,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m101011_0	),
Adb40101111100	(	adb40101111100,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m101011_0	),
Adb40101111101	(	adb40101111101,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m101011_0	),
Adb40101111110	(	adb40101111110,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m101011_0	),
Adb40101111111	(	adb40101111111,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m101011_0	),
Adb40110000000	(	adb40110000000,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m100011_0	),
Adb40110000001	(	adb40110000001,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m100011_0	),
Adb40110000010	(	adb40110000010,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m100011_0	),
Adb40110000011	(	adb40110000011,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m100011_0	),
Adb40110000100	(	adb40110000100,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m100011_0	),
Adb40110000101	(	adb40110000101,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m100011_0	),
Adb40110000110	(	adb40110000110,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m100011_0	),
Adb40110000111	(	adb40110000111,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m100011_0	),
Adb40110001000	(	adb40110001000,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m100011_0	),
Adb40110001001	(	adb40110001001,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m100011_0	),
Adb40110001010	(	adb40110001010,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m100011_0	),
Adb40110001011	(	adb40110001011,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m100011_0	),
Adb40110001100	(	adb40110001100,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m100011_0	),
Adb40110001101	(	adb40110001101,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m100011_0	),
Adb40110001110	(	adb40110001110,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m100011_0	),
Adb40110001111	(	adb40110001111,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m100011_0	),
Adb40110010000	(	adb40110010000,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m100011_0	),
Adb40110010001	(	adb40110010001,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m100011_0	),
Adb40110010010	(	adb40110010010,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m100011_0	),
Adb40110010011	(	adb40110010011,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m100011_0	),
Adb40110010100	(	adb40110010100,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m100011_0	),
Adb40110010101	(	adb40110010101,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m100011_0	),
Adb40110010110	(	adb40110010110,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m100011_0	),
Adb40110010111	(	adb40110010111,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m100011_0	),
Adb40110011000	(	adb40110011000,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m100011_0	),
Adb40110011001	(	adb40110011001,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m100011_0	),
Adb40110011010	(	adb40110011010,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m100011_0	),
Adb40110011011	(	adb40110011011,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m100011_0	),
Adb40110011100	(	adb40110011100,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m100011_0	),
Adb40110011101	(	adb40110011101,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m100011_0	),
Adb40110011110	(	adb40110011110,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m100011_0	),
Adb40110011111	(	adb40110011111,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m100011_0	),
Adb40110100000	(	adb40110100000,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m100011_0	),
Adb40110100001	(	adb40110100001,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m100011_0	),
Adb40110100010	(	adb40110100010,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m100011_0	),
Adb40110100011	(	adb40110100011,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m100011_0	),
Adb40110100100	(	adb40110100100,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m100011_0	),
Adb40110100101	(	adb40110100101,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m100011_0	),
Adb40110100110	(	adb40110100110,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m100011_0	),
Adb40110100111	(	adb40110100111,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m100011_0	),
Adb40110101000	(	adb40110101000,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m100011_0	),
Adb40110101001	(	adb40110101001,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m100011_0	),
Adb40110101010	(	adb40110101010,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m100011_0	),
Adb40110101011	(	adb40110101011,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m100011_0	),
Adb40110101100	(	adb40110101100,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m100011_0	),
Adb40110101101	(	adb40110101101,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m100011_0	),
Adb40110101110	(	adb40110101110,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m100011_0	),
Adb40110101111	(	adb40110101111,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m100011_0	),
Adb40110110000	(	adb40110110000,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m100011_0	),
Adb40110110001	(	adb40110110001,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m100011_0	),
Adb40110110010	(	adb40110110010,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m100011_0	),
Adb40110110011	(	adb40110110011,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m100011_0	),
Adb40110110100	(	adb40110110100,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m100011_0	),
Adb40110110101	(	adb40110110101,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m100011_0	),
Adb40110110110	(	adb40110110110,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m100011_0	),
Adb40110110111	(	adb40110110111,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m100011_0	),
Adb40110111000	(	adb40110111000,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m100011_0	),
Adb40110111001	(	adb40110111001,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m100011_0	),
Adb40110111010	(	adb40110111010,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m100011_0	),
Adb40110111011	(	adb40110111011,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m100011_0	),
Adb40110111100	(	adb40110111100,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m100011_0	),
Adb40110111101	(	adb40110111101,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m100011_0	),
Adb40110111110	(	adb40110111110,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m100011_0	),
Adb40110111111	(	adb40110111111,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m100011_0	),
Adb40111000000	(	adb40111000000,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m100011_0	),
Adb40111000001	(	adb40111000001,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m100011_0	),
Adb40111000010	(	adb40111000010,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m100011_0	),
Adb40111000011	(	adb40111000011,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m100011_0	),
Adb40111000100	(	adb40111000100,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m100011_0	),
Adb40111000101	(	adb40111000101,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m100011_0	),
Adb40111000110	(	adb40111000110,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m100011_0	),
Adb40111000111	(	adb40111000111,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m100011_0	),
Adb40111001000	(	adb40111001000,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m100011_0	),
Adb40111001001	(	adb40111001001,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m100011_0	),
Adb40111001010	(	adb40111001010,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m100011_0	),
Adb40111001011	(	adb40111001011,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m100011_0	),
Adb40111001100	(	adb40111001100,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m100011_0	),
Adb40111001101	(	adb40111001101,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m100011_0	),
Adb40111001110	(	adb40111001110,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m100011_0	),
Adb40111001111	(	adb40111001111,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m100011_0	),
Adb40111010000	(	adb40111010000,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m100011_0	),
Adb40111010001	(	adb40111010001,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m100011_0	),
Adb40111010010	(	adb40111010010,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m100011_0	),
Adb40111010011	(	adb40111010011,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m100011_0	),
Adb40111010100	(	adb40111010100,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m100011_0	),
Adb40111010101	(	adb40111010101,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m100011_0	),
Adb40111010110	(	adb40111010110,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m100011_0	),
Adb40111010111	(	adb40111010111,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m100011_0	),
Adb40111011000	(	adb40111011000,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m100011_0	),
Adb40111011001	(	adb40111011001,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m100011_0	),
Adb40111011010	(	adb40111011010,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m100011_0	),
Adb40111011011	(	adb40111011011,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m100011_0	),
Adb40111011100	(	adb40111011100,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m100011_0	),
Adb40111011101	(	adb40111011101,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m100011_0	),
Adb40111011110	(	adb40111011110,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m100011_0	),
Adb40111011111	(	adb40111011111,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m100011_0	),
Adb40111100000	(	adb40111100000,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m100011_0	),
Adb40111100001	(	adb40111100001,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m100011_0	),
Adb40111100010	(	adb40111100010,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m100011_0	),
Adb40111100011	(	adb40111100011,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m100011_0	),
Adb40111100100	(	adb40111100100,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m100011_0	),
Adb40111100101	(	adb40111100101,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m100011_0	),
Adb40111100110	(	adb40111100110,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m100011_0	),
Adb40111100111	(	adb40111100111,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m100011_0	),
Adb40111101000	(	adb40111101000,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m100011_0	),
Adb40111101001	(	adb40111101001,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m100011_0	),
Adb40111101010	(	adb40111101010,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m100011_0	),
Adb40111101011	(	adb40111101011,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m100011_0	),
Adb40111101100	(	adb40111101100,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m100011_0	),
Adb40111101101	(	adb40111101101,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m100011_0	),
Adb40111101110	(	adb40111101110,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m100011_0	),
Adb40111101111	(	adb40111101111,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m100011_0	),
Adb40111110000	(	adb40111110000,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m100011_0	),
Adb40111110001	(	adb40111110001,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m100011_0	),
Adb40111110010	(	adb40111110010,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m100011_0	),
Adb40111110011	(	adb40111110011,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m100011_0	),
Adb40111110100	(	adb40111110100,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m100011_0	),
Adb40111110101	(	adb40111110101,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m100011_0	),
Adb40111110110	(	adb40111110110,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m100011_0	),
Adb40111110111	(	adb40111110111,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m100011_0	),
Adb40111111000	(	adb40111111000,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m100011_0	),
Adb40111111001	(	adb40111111001,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m100011_0	),
Adb40111111010	(	adb40111111010,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m100011_0	),
Adb40111111011	(	adb40111111011,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m100011_0	),
Adb40111111100	(	adb40111111100,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m100011_0	),
Adb40111111101	(	adb40111111101,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m100011_0	),
Adb40111111110	(	adb40111111110,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m100011_0	),
Adb40111111111	(	adb40111111111,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m100011_0	),
Adb41000000000	(	adb41000000000,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m011011_0	),
Adb41000000001	(	adb41000000001,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m011011_0	),
Adb41000000010	(	adb41000000010,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m011011_0	),
Adb41000000011	(	adb41000000011,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m011011_0	),
Adb41000000100	(	adb41000000100,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m011011_0	),
Adb41000000101	(	adb41000000101,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m011011_0	),
Adb41000000110	(	adb41000000110,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m011011_0	),
Adb41000000111	(	adb41000000111,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m011011_0	),
Adb41000001000	(	adb41000001000,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m011011_0	),
Adb41000001001	(	adb41000001001,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m011011_0	),
Adb41000001010	(	adb41000001010,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m011011_0	),
Adb41000001011	(	adb41000001011,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m011011_0	),
Adb41000001100	(	adb41000001100,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m011011_0	),
Adb41000001101	(	adb41000001101,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m011011_0	),
Adb41000001110	(	adb41000001110,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m011011_0	),
Adb41000001111	(	adb41000001111,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m011011_0	),
Adb41000010000	(	adb41000010000,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m011011_0	),
Adb41000010001	(	adb41000010001,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m011011_0	),
Adb41000010010	(	adb41000010010,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m011011_0	),
Adb41000010011	(	adb41000010011,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m011011_0	),
Adb41000010100	(	adb41000010100,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m011011_0	),
Adb41000010101	(	adb41000010101,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m011011_0	),
Adb41000010110	(	adb41000010110,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m011011_0	),
Adb41000010111	(	adb41000010111,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m011011_0	),
Adb41000011000	(	adb41000011000,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m011011_0	),
Adb41000011001	(	adb41000011001,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m011011_0	),
Adb41000011010	(	adb41000011010,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m011011_0	),
Adb41000011011	(	adb41000011011,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m011011_0	),
Adb41000011100	(	adb41000011100,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m011011_0	),
Adb41000011101	(	adb41000011101,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m011011_0	),
Adb41000011110	(	adb41000011110,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m011011_0	),
Adb41000011111	(	adb41000011111,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m011011_0	),
Adb41000100000	(	adb41000100000,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m011011_0	),
Adb41000100001	(	adb41000100001,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m011011_0	),
Adb41000100010	(	adb41000100010,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m011011_0	),
Adb41000100011	(	adb41000100011,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m011011_0	),
Adb41000100100	(	adb41000100100,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m011011_0	),
Adb41000100101	(	adb41000100101,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m011011_0	),
Adb41000100110	(	adb41000100110,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m011011_0	),
Adb41000100111	(	adb41000100111,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m011011_0	),
Adb41000101000	(	adb41000101000,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m011011_0	),
Adb41000101001	(	adb41000101001,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m011011_0	),
Adb41000101010	(	adb41000101010,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m011011_0	),
Adb41000101011	(	adb41000101011,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m011011_0	),
Adb41000101100	(	adb41000101100,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m011011_0	),
Adb41000101101	(	adb41000101101,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m011011_0	),
Adb41000101110	(	adb41000101110,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m011011_0	),
Adb41000101111	(	adb41000101111,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m011011_0	),
Adb41000110000	(	adb41000110000,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m011011_0	),
Adb41000110001	(	adb41000110001,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m011011_0	),
Adb41000110010	(	adb41000110010,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m011011_0	),
Adb41000110011	(	adb41000110011,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m011011_0	),
Adb41000110100	(	adb41000110100,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m011011_0	),
Adb41000110101	(	adb41000110101,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m011011_0	),
Adb41000110110	(	adb41000110110,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m011011_0	),
Adb41000110111	(	adb41000110111,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m011011_0	),
Adb41000111000	(	adb41000111000,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m011011_0	),
Adb41000111001	(	adb41000111001,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m011011_0	),
Adb41000111010	(	adb41000111010,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m011011_0	),
Adb41000111011	(	adb41000111011,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m011011_0	),
Adb41000111100	(	adb41000111100,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m011011_0	),
Adb41000111101	(	adb41000111101,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m011011_0	),
Adb41000111110	(	adb41000111110,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m011011_0	),
Adb41000111111	(	adb41000111111,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m011011_0	),
Adb41001000000	(	adb41001000000,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m011011_0	),
Adb41001000001	(	adb41001000001,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m011011_0	),
Adb41001000010	(	adb41001000010,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m011011_0	),
Adb41001000011	(	adb41001000011,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m011011_0	),
Adb41001000100	(	adb41001000100,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m011011_0	),
Adb41001000101	(	adb41001000101,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m011011_0	),
Adb41001000110	(	adb41001000110,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m011011_0	),
Adb41001000111	(	adb41001000111,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m011011_0	),
Adb41001001000	(	adb41001001000,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m011011_0	),
Adb41001001001	(	adb41001001001,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m011011_0	),
Adb41001001010	(	adb41001001010,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m011011_0	),
Adb41001001011	(	adb41001001011,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m011011_0	),
Adb41001001100	(	adb41001001100,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m011011_0	),
Adb41001001101	(	adb41001001101,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m011011_0	),
Adb41001001110	(	adb41001001110,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m011011_0	),
Adb41001001111	(	adb41001001111,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m011011_0	),
Adb41001010000	(	adb41001010000,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m011011_0	),
Adb41001010001	(	adb41001010001,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m011011_0	),
Adb41001010010	(	adb41001010010,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m011011_0	),
Adb41001010011	(	adb41001010011,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m011011_0	),
Adb41001010100	(	adb41001010100,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m011011_0	),
Adb41001010101	(	adb41001010101,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m011011_0	),
Adb41001010110	(	adb41001010110,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m011011_0	),
Adb41001010111	(	adb41001010111,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m011011_0	),
Adb41001011000	(	adb41001011000,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m011011_0	),
Adb41001011001	(	adb41001011001,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m011011_0	),
Adb41001011010	(	adb41001011010,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m011011_0	),
Adb41001011011	(	adb41001011011,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m011011_0	),
Adb41001011100	(	adb41001011100,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m011011_0	),
Adb41001011101	(	adb41001011101,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m011011_0	),
Adb41001011110	(	adb41001011110,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m011011_0	),
Adb41001011111	(	adb41001011111,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m011011_0	),
Adb41001100000	(	adb41001100000,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m011011_0	),
Adb41001100001	(	adb41001100001,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m011011_0	),
Adb41001100010	(	adb41001100010,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m011011_0	),
Adb41001100011	(	adb41001100011,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m011011_0	),
Adb41001100100	(	adb41001100100,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m011011_0	),
Adb41001100101	(	adb41001100101,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m011011_0	),
Adb41001100110	(	adb41001100110,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m011011_0	),
Adb41001100111	(	adb41001100111,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m011011_0	),
Adb41001101000	(	adb41001101000,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m011011_0	),
Adb41001101001	(	adb41001101001,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m011011_0	),
Adb41001101010	(	adb41001101010,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m011011_0	),
Adb41001101011	(	adb41001101011,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m011011_0	),
Adb41001101100	(	adb41001101100,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m011011_0	),
Adb41001101101	(	adb41001101101,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m011011_0	),
Adb41001101110	(	adb41001101110,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m011011_0	),
Adb41001101111	(	adb41001101111,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m011011_0	),
Adb41001110000	(	adb41001110000,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m011011_0	),
Adb41001110001	(	adb41001110001,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m011011_0	),
Adb41001110010	(	adb41001110010,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m011011_0	),
Adb41001110011	(	adb41001110011,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m011011_0	),
Adb41001110100	(	adb41001110100,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m011011_0	),
Adb41001110101	(	adb41001110101,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m011011_0	),
Adb41001110110	(	adb41001110110,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m011011_0	),
Adb41001110111	(	adb41001110111,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m011011_0	),
Adb41001111000	(	adb41001111000,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m011011_0	),
Adb41001111001	(	adb41001111001,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m011011_0	),
Adb41001111010	(	adb41001111010,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m011011_0	),
Adb41001111011	(	adb41001111011,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m011011_0	),
Adb41001111100	(	adb41001111100,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m011011_0	),
Adb41001111101	(	adb41001111101,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m011011_0	),
Adb41001111110	(	adb41001111110,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m011011_0	),
Adb41001111111	(	adb41001111111,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m011011_0	),
Adb41010000000	(	adb41010000000,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m010011_0	),
Adb41010000001	(	adb41010000001,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m010011_0	),
Adb41010000010	(	adb41010000010,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m010011_0	),
Adb41010000011	(	adb41010000011,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m010011_0	),
Adb41010000100	(	adb41010000100,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m010011_0	),
Adb41010000101	(	adb41010000101,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m010011_0	),
Adb41010000110	(	adb41010000110,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m010011_0	),
Adb41010000111	(	adb41010000111,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m010011_0	),
Adb41010001000	(	adb41010001000,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m010011_0	),
Adb41010001001	(	adb41010001001,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m010011_0	),
Adb41010001010	(	adb41010001010,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m010011_0	),
Adb41010001011	(	adb41010001011,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m010011_0	),
Adb41010001100	(	adb41010001100,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m010011_0	),
Adb41010001101	(	adb41010001101,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m010011_0	),
Adb41010001110	(	adb41010001110,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m010011_0	),
Adb41010001111	(	adb41010001111,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m010011_0	),
Adb41010010000	(	adb41010010000,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m010011_0	),
Adb41010010001	(	adb41010010001,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m010011_0	),
Adb41010010010	(	adb41010010010,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m010011_0	),
Adb41010010011	(	adb41010010011,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m010011_0	),
Adb41010010100	(	adb41010010100,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m010011_0	),
Adb41010010101	(	adb41010010101,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m010011_0	),
Adb41010010110	(	adb41010010110,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m010011_0	),
Adb41010010111	(	adb41010010111,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m010011_0	),
Adb41010011000	(	adb41010011000,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m010011_0	),
Adb41010011001	(	adb41010011001,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m010011_0	),
Adb41010011010	(	adb41010011010,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m010011_0	),
Adb41010011011	(	adb41010011011,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m010011_0	),
Adb41010011100	(	adb41010011100,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m010011_0	),
Adb41010011101	(	adb41010011101,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m010011_0	),
Adb41010011110	(	adb41010011110,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m010011_0	),
Adb41010011111	(	adb41010011111,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m010011_0	),
Adb41010100000	(	adb41010100000,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m010011_0	),
Adb41010100001	(	adb41010100001,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m010011_0	),
Adb41010100010	(	adb41010100010,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m010011_0	),
Adb41010100011	(	adb41010100011,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m010011_0	),
Adb41010100100	(	adb41010100100,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m010011_0	),
Adb41010100101	(	adb41010100101,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m010011_0	),
Adb41010100110	(	adb41010100110,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m010011_0	),
Adb41010100111	(	adb41010100111,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m010011_0	),
Adb41010101000	(	adb41010101000,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m010011_0	),
Adb41010101001	(	adb41010101001,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m010011_0	),
Adb41010101010	(	adb41010101010,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m010011_0	),
Adb41010101011	(	adb41010101011,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m010011_0	),
Adb41010101100	(	adb41010101100,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m010011_0	),
Adb41010101101	(	adb41010101101,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m010011_0	),
Adb41010101110	(	adb41010101110,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m010011_0	),
Adb41010101111	(	adb41010101111,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m010011_0	),
Adb41010110000	(	adb41010110000,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m010011_0	),
Adb41010110001	(	adb41010110001,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m010011_0	),
Adb41010110010	(	adb41010110010,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m010011_0	),
Adb41010110011	(	adb41010110011,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m010011_0	),
Adb41010110100	(	adb41010110100,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m010011_0	),
Adb41010110101	(	adb41010110101,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m010011_0	),
Adb41010110110	(	adb41010110110,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m010011_0	),
Adb41010110111	(	adb41010110111,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m010011_0	),
Adb41010111000	(	adb41010111000,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m010011_0	),
Adb41010111001	(	adb41010111001,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m010011_0	),
Adb41010111010	(	adb41010111010,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m010011_0	),
Adb41010111011	(	adb41010111011,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m010011_0	),
Adb41010111100	(	adb41010111100,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m010011_0	),
Adb41010111101	(	adb41010111101,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m010011_0	),
Adb41010111110	(	adb41010111110,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m010011_0	),
Adb41010111111	(	adb41010111111,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m010011_0	),
Adb41011000000	(	adb41011000000,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m010011_0	),
Adb41011000001	(	adb41011000001,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m010011_0	),
Adb41011000010	(	adb41011000010,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m010011_0	),
Adb41011000011	(	adb41011000011,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m010011_0	),
Adb41011000100	(	adb41011000100,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m010011_0	),
Adb41011000101	(	adb41011000101,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m010011_0	),
Adb41011000110	(	adb41011000110,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m010011_0	),
Adb41011000111	(	adb41011000111,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m010011_0	),
Adb41011001000	(	adb41011001000,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m010011_0	),
Adb41011001001	(	adb41011001001,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m010011_0	),
Adb41011001010	(	adb41011001010,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m010011_0	),
Adb41011001011	(	adb41011001011,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m010011_0	),
Adb41011001100	(	adb41011001100,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m010011_0	),
Adb41011001101	(	adb41011001101,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m010011_0	),
Adb41011001110	(	adb41011001110,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m010011_0	),
Adb41011001111	(	adb41011001111,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m010011_0	),
Adb41011010000	(	adb41011010000,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m010011_0	),
Adb41011010001	(	adb41011010001,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m010011_0	),
Adb41011010010	(	adb41011010010,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m010011_0	),
Adb41011010011	(	adb41011010011,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m010011_0	),
Adb41011010100	(	adb41011010100,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m010011_0	),
Adb41011010101	(	adb41011010101,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m010011_0	),
Adb41011010110	(	adb41011010110,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m010011_0	),
Adb41011010111	(	adb41011010111,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m010011_0	),
Adb41011011000	(	adb41011011000,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m010011_0	),
Adb41011011001	(	adb41011011001,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m010011_0	),
Adb41011011010	(	adb41011011010,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m010011_0	),
Adb41011011011	(	adb41011011011,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m010011_0	),
Adb41011011100	(	adb41011011100,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m010011_0	),
Adb41011011101	(	adb41011011101,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m010011_0	),
Adb41011011110	(	adb41011011110,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m010011_0	),
Adb41011011111	(	adb41011011111,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m010011_0	),
Adb41011100000	(	adb41011100000,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m010011_0	),
Adb41011100001	(	adb41011100001,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m010011_0	),
Adb41011100010	(	adb41011100010,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m010011_0	),
Adb41011100011	(	adb41011100011,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m010011_0	),
Adb41011100100	(	adb41011100100,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m010011_0	),
Adb41011100101	(	adb41011100101,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m010011_0	),
Adb41011100110	(	adb41011100110,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m010011_0	),
Adb41011100111	(	adb41011100111,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m010011_0	),
Adb41011101000	(	adb41011101000,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m010011_0	),
Adb41011101001	(	adb41011101001,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m010011_0	),
Adb41011101010	(	adb41011101010,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m010011_0	),
Adb41011101011	(	adb41011101011,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m010011_0	),
Adb41011101100	(	adb41011101100,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m010011_0	),
Adb41011101101	(	adb41011101101,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m010011_0	),
Adb41011101110	(	adb41011101110,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m010011_0	),
Adb41011101111	(	adb41011101111,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m010011_0	),
Adb41011110000	(	adb41011110000,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m010011_0	),
Adb41011110001	(	adb41011110001,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m010011_0	),
Adb41011110010	(	adb41011110010,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m010011_0	),
Adb41011110011	(	adb41011110011,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m010011_0	),
Adb41011110100	(	adb41011110100,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m010011_0	),
Adb41011110101	(	adb41011110101,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m010011_0	),
Adb41011110110	(	adb41011110110,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m010011_0	),
Adb41011110111	(	adb41011110111,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m010011_0	),
Adb41011111000	(	adb41011111000,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m010011_0	),
Adb41011111001	(	adb41011111001,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m010011_0	),
Adb41011111010	(	adb41011111010,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m010011_0	),
Adb41011111011	(	adb41011111011,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m010011_0	),
Adb41011111100	(	adb41011111100,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m010011_0	),
Adb41011111101	(	adb41011111101,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m010011_0	),
Adb41011111110	(	adb41011111110,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m010011_0	),
Adb41011111111	(	adb41011111111,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m010011_0	),
Adb41100000000	(	adb41100000000,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m001011_0	),
Adb41100000001	(	adb41100000001,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m001011_0	),
Adb41100000010	(	adb41100000010,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m001011_0	),
Adb41100000011	(	adb41100000011,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m001011_0	),
Adb41100000100	(	adb41100000100,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m001011_0	),
Adb41100000101	(	adb41100000101,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m001011_0	),
Adb41100000110	(	adb41100000110,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m001011_0	),
Adb41100000111	(	adb41100000111,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m001011_0	),
Adb41100001000	(	adb41100001000,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m001011_0	),
Adb41100001001	(	adb41100001001,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m001011_0	),
Adb41100001010	(	adb41100001010,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m001011_0	),
Adb41100001011	(	adb41100001011,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m001011_0	),
Adb41100001100	(	adb41100001100,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m001011_0	),
Adb41100001101	(	adb41100001101,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m001011_0	),
Adb41100001110	(	adb41100001110,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m001011_0	),
Adb41100001111	(	adb41100001111,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m001011_0	),
Adb41100010000	(	adb41100010000,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m001011_0	),
Adb41100010001	(	adb41100010001,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m001011_0	),
Adb41100010010	(	adb41100010010,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m001011_0	),
Adb41100010011	(	adb41100010011,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m001011_0	),
Adb41100010100	(	adb41100010100,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m001011_0	),
Adb41100010101	(	adb41100010101,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m001011_0	),
Adb41100010110	(	adb41100010110,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m001011_0	),
Adb41100010111	(	adb41100010111,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m001011_0	),
Adb41100011000	(	adb41100011000,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m001011_0	),
Adb41100011001	(	adb41100011001,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m001011_0	),
Adb41100011010	(	adb41100011010,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m001011_0	),
Adb41100011011	(	adb41100011011,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m001011_0	),
Adb41100011100	(	adb41100011100,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m001011_0	),
Adb41100011101	(	adb41100011101,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m001011_0	),
Adb41100011110	(	adb41100011110,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m001011_0	),
Adb41100011111	(	adb41100011111,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m001011_0	),
Adb41100100000	(	adb41100100000,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m001011_0	),
Adb41100100001	(	adb41100100001,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m001011_0	),
Adb41100100010	(	adb41100100010,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m001011_0	),
Adb41100100011	(	adb41100100011,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m001011_0	),
Adb41100100100	(	adb41100100100,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m001011_0	),
Adb41100100101	(	adb41100100101,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m001011_0	),
Adb41100100110	(	adb41100100110,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m001011_0	),
Adb41100100111	(	adb41100100111,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m001011_0	),
Adb41100101000	(	adb41100101000,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m001011_0	),
Adb41100101001	(	adb41100101001,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m001011_0	),
Adb41100101010	(	adb41100101010,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m001011_0	),
Adb41100101011	(	adb41100101011,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m001011_0	),
Adb41100101100	(	adb41100101100,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m001011_0	),
Adb41100101101	(	adb41100101101,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m001011_0	),
Adb41100101110	(	adb41100101110,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m001011_0	),
Adb41100101111	(	adb41100101111,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m001011_0	),
Adb41100110000	(	adb41100110000,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m001011_0	),
Adb41100110001	(	adb41100110001,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m001011_0	),
Adb41100110010	(	adb41100110010,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m001011_0	),
Adb41100110011	(	adb41100110011,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m001011_0	),
Adb41100110100	(	adb41100110100,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m001011_0	),
Adb41100110101	(	adb41100110101,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m001011_0	),
Adb41100110110	(	adb41100110110,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m001011_0	),
Adb41100110111	(	adb41100110111,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m001011_0	),
Adb41100111000	(	adb41100111000,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m001011_0	),
Adb41100111001	(	adb41100111001,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m001011_0	),
Adb41100111010	(	adb41100111010,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m001011_0	),
Adb41100111011	(	adb41100111011,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m001011_0	),
Adb41100111100	(	adb41100111100,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m001011_0	),
Adb41100111101	(	adb41100111101,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m001011_0	),
Adb41100111110	(	adb41100111110,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m001011_0	),
Adb41100111111	(	adb41100111111,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m001011_0	),
Adb41101000000	(	adb41101000000,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m001011_0	),
Adb41101000001	(	adb41101000001,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m001011_0	),
Adb41101000010	(	adb41101000010,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m001011_0	),
Adb41101000011	(	adb41101000011,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m001011_0	),
Adb41101000100	(	adb41101000100,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m001011_0	),
Adb41101000101	(	adb41101000101,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m001011_0	),
Adb41101000110	(	adb41101000110,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m001011_0	),
Adb41101000111	(	adb41101000111,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m001011_0	),
Adb41101001000	(	adb41101001000,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m001011_0	),
Adb41101001001	(	adb41101001001,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m001011_0	),
Adb41101001010	(	adb41101001010,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m001011_0	),
Adb41101001011	(	adb41101001011,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m001011_0	),
Adb41101001100	(	adb41101001100,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m001011_0	),
Adb41101001101	(	adb41101001101,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m001011_0	),
Adb41101001110	(	adb41101001110,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m001011_0	),
Adb41101001111	(	adb41101001111,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m001011_0	),
Adb41101010000	(	adb41101010000,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m001011_0	),
Adb41101010001	(	adb41101010001,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m001011_0	),
Adb41101010010	(	adb41101010010,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m001011_0	),
Adb41101010011	(	adb41101010011,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m001011_0	),
Adb41101010100	(	adb41101010100,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m001011_0	),
Adb41101010101	(	adb41101010101,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m001011_0	),
Adb41101010110	(	adb41101010110,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m001011_0	),
Adb41101010111	(	adb41101010111,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m001011_0	),
Adb41101011000	(	adb41101011000,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m001011_0	),
Adb41101011001	(	adb41101011001,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m001011_0	),
Adb41101011010	(	adb41101011010,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m001011_0	),
Adb41101011011	(	adb41101011011,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m001011_0	),
Adb41101011100	(	adb41101011100,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m001011_0	),
Adb41101011101	(	adb41101011101,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m001011_0	),
Adb41101011110	(	adb41101011110,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m001011_0	),
Adb41101011111	(	adb41101011111,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m001011_0	),
Adb41101100000	(	adb41101100000,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m001011_0	),
Adb41101100001	(	adb41101100001,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m001011_0	),
Adb41101100010	(	adb41101100010,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m001011_0	),
Adb41101100011	(	adb41101100011,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m001011_0	),
Adb41101100100	(	adb41101100100,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m001011_0	),
Adb41101100101	(	adb41101100101,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m001011_0	),
Adb41101100110	(	adb41101100110,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m001011_0	),
Adb41101100111	(	adb41101100111,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m001011_0	),
Adb41101101000	(	adb41101101000,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m001011_0	),
Adb41101101001	(	adb41101101001,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m001011_0	),
Adb41101101010	(	adb41101101010,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m001011_0	),
Adb41101101011	(	adb41101101011,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m001011_0	),
Adb41101101100	(	adb41101101100,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m001011_0	),
Adb41101101101	(	adb41101101101,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m001011_0	),
Adb41101101110	(	adb41101101110,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m001011_0	),
Adb41101101111	(	adb41101101111,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m001011_0	),
Adb41101110000	(	adb41101110000,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m001011_0	),
Adb41101110001	(	adb41101110001,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m001011_0	),
Adb41101110010	(	adb41101110010,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m001011_0	),
Adb41101110011	(	adb41101110011,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m001011_0	),
Adb41101110100	(	adb41101110100,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m001011_0	),
Adb41101110101	(	adb41101110101,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m001011_0	),
Adb41101110110	(	adb41101110110,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m001011_0	),
Adb41101110111	(	adb41101110111,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m001011_0	),
Adb41101111000	(	adb41101111000,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m001011_0	),
Adb41101111001	(	adb41101111001,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m001011_0	),
Adb41101111010	(	adb41101111010,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m001011_0	),
Adb41101111011	(	adb41101111011,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m001011_0	),
Adb41101111100	(	adb41101111100,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m001011_0	),
Adb41101111101	(	adb41101111101,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m001011_0	),
Adb41101111110	(	adb41101111110,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m001011_0	),
Adb41101111111	(	adb41101111111,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m001011_0	),
Adb41110000000	(	adb41110000000,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m000011_0	),
Adb41110000001	(	adb41110000001,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m000011_0	),
Adb41110000010	(	adb41110000010,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m000011_0	),
Adb41110000011	(	adb41110000011,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m000011_0	),
Adb41110000100	(	adb41110000100,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m000011_0	),
Adb41110000101	(	adb41110000101,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m000011_0	),
Adb41110000110	(	adb41110000110,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m000011_0	),
Adb41110000111	(	adb41110000111,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m000011_0	),
Adb41110001000	(	adb41110001000,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m000011_0	),
Adb41110001001	(	adb41110001001,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m000011_0	),
Adb41110001010	(	adb41110001010,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m000011_0	),
Adb41110001011	(	adb41110001011,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m000011_0	),
Adb41110001100	(	adb41110001100,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m000011_0	),
Adb41110001101	(	adb41110001101,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m000011_0	),
Adb41110001110	(	adb41110001110,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m000011_0	),
Adb41110001111	(	adb41110001111,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m000011_0	),
Adb41110010000	(	adb41110010000,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m000011_0	),
Adb41110010001	(	adb41110010001,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m000011_0	),
Adb41110010010	(	adb41110010010,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m000011_0	),
Adb41110010011	(	adb41110010011,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m000011_0	),
Adb41110010100	(	adb41110010100,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m000011_0	),
Adb41110010101	(	adb41110010101,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m000011_0	),
Adb41110010110	(	adb41110010110,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m000011_0	),
Adb41110010111	(	adb41110010111,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m000011_0	),
Adb41110011000	(	adb41110011000,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m000011_0	),
Adb41110011001	(	adb41110011001,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m000011_0	),
Adb41110011010	(	adb41110011010,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m000011_0	),
Adb41110011011	(	adb41110011011,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m000011_0	),
Adb41110011100	(	adb41110011100,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m000011_0	),
Adb41110011101	(	adb41110011101,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m000011_0	),
Adb41110011110	(	adb41110011110,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m000011_0	),
Adb41110011111	(	adb41110011111,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m000011_0	),
Adb41110100000	(	adb41110100000,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m000011_0	),
Adb41110100001	(	adb41110100001,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m000011_0	),
Adb41110100010	(	adb41110100010,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m000011_0	),
Adb41110100011	(	adb41110100011,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m000011_0	),
Adb41110100100	(	adb41110100100,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m000011_0	),
Adb41110100101	(	adb41110100101,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m000011_0	),
Adb41110100110	(	adb41110100110,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m000011_0	),
Adb41110100111	(	adb41110100111,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m000011_0	),
Adb41110101000	(	adb41110101000,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m000011_0	),
Adb41110101001	(	adb41110101001,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m000011_0	),
Adb41110101010	(	adb41110101010,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m000011_0	),
Adb41110101011	(	adb41110101011,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m000011_0	),
Adb41110101100	(	adb41110101100,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m000011_0	),
Adb41110101101	(	adb41110101101,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m000011_0	),
Adb41110101110	(	adb41110101110,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m000011_0	),
Adb41110101111	(	adb41110101111,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m000011_0	),
Adb41110110000	(	adb41110110000,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m000011_0	),
Adb41110110001	(	adb41110110001,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m000011_0	),
Adb41110110010	(	adb41110110010,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m000011_0	),
Adb41110110011	(	adb41110110011,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m000011_0	),
Adb41110110100	(	adb41110110100,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m000011_0	),
Adb41110110101	(	adb41110110101,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m000011_0	),
Adb41110110110	(	adb41110110110,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m000011_0	),
Adb41110110111	(	adb41110110111,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m000011_0	),
Adb41110111000	(	adb41110111000,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m000011_0	),
Adb41110111001	(	adb41110111001,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m000011_0	),
Adb41110111010	(	adb41110111010,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m000011_0	),
Adb41110111011	(	adb41110111011,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m000011_0	),
Adb41110111100	(	adb41110111100,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m000011_0	),
Adb41110111101	(	adb41110111101,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m000011_0	),
Adb41110111110	(	adb41110111110,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m000011_0	),
Adb41110111111	(	adb41110111111,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m000011_0	),
Adb41111000000	(	adb41111000000,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m000011_0	),
Adb41111000001	(	adb41111000001,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m000011_0	),
Adb41111000010	(	adb41111000010,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m000011_0	),
Adb41111000011	(	adb41111000011,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m000011_0	),
Adb41111000100	(	adb41111000100,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m000011_0	),
Adb41111000101	(	adb41111000101,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m000011_0	),
Adb41111000110	(	adb41111000110,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m000011_0	),
Adb41111000111	(	adb41111000111,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m000011_0	),
Adb41111001000	(	adb41111001000,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m000011_0	),
Adb41111001001	(	adb41111001001,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m000011_0	),
Adb41111001010	(	adb41111001010,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m000011_0	),
Adb41111001011	(	adb41111001011,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m000011_0	),
Adb41111001100	(	adb41111001100,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m000011_0	),
Adb41111001101	(	adb41111001101,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m000011_0	),
Adb41111001110	(	adb41111001110,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m000011_0	),
Adb41111001111	(	adb41111001111,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m000011_0	),
Adb41111010000	(	adb41111010000,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m000011_0	),
Adb41111010001	(	adb41111010001,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m000011_0	),
Adb41111010010	(	adb41111010010,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m000011_0	),
Adb41111010011	(	adb41111010011,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m000011_0	),
Adb41111010100	(	adb41111010100,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m000011_0	),
Adb41111010101	(	adb41111010101,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m000011_0	),
Adb41111010110	(	adb41111010110,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m000011_0	),
Adb41111010111	(	adb41111010111,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m000011_0	),
Adb41111011000	(	adb41111011000,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m000011_0	),
Adb41111011001	(	adb41111011001,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m000011_0	),
Adb41111011010	(	adb41111011010,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m000011_0	),
Adb41111011011	(	adb41111011011,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m000011_0	),
Adb41111011100	(	adb41111011100,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m000011_0	),
Adb41111011101	(	adb41111011101,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m000011_0	),
Adb41111011110	(	adb41111011110,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m000011_0	),
Adb41111011111	(	adb41111011111,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m000011_0	),
Adb41111100000	(	adb41111100000,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m000011_0	),
Adb41111100001	(	adb41111100001,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m000011_0	),
Adb41111100010	(	adb41111100010,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m000011_0	),
Adb41111100011	(	adb41111100011,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m000011_0	),
Adb41111100100	(	adb41111100100,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m000011_0	),
Adb41111100101	(	adb41111100101,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m000011_0	),
Adb41111100110	(	adb41111100110,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m000011_0	),
Adb41111100111	(	adb41111100111,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m000011_0	),
Adb41111101000	(	adb41111101000,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m000011_0	),
Adb41111101001	(	adb41111101001,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m000011_0	),
Adb41111101010	(	adb41111101010,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m000011_0	),
Adb41111101011	(	adb41111101011,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m000011_0	),
Adb41111101100	(	adb41111101100,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m000011_0	),
Adb41111101101	(	adb41111101101,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m000011_0	),
Adb41111101110	(	adb41111101110,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m000011_0	),
Adb41111101111	(	adb41111101111,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m000011_0	),
Adb41111110000	(	adb41111110000,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m000011_0	),
Adb41111110001	(	adb41111110001,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m000011_0	),
Adb41111110010	(	adb41111110010,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m000011_0	),
Adb41111110011	(	adb41111110011,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m000011_0	),
Adb41111110100	(	adb41111110100,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m000011_0	),
Adb41111110101	(	adb41111110101,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m000011_0	),
Adb41111110110	(	adb41111110110,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m000011_0	),
Adb41111110111	(	adb41111110111,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m000011_0	),
Adb41111111000	(	adb41111111000,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m000011_0	),
Adb41111111001	(	adb41111111001,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m000011_0	),
Adb41111111010	(	adb41111111010,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m000011_0	),
Adb41111111011	(	adb41111111011,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m000011_0	),
Adb41111111100	(	adb41111111100,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m000011_0	),
Adb41111111101	(	adb41111111101,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m000011_0	),
Adb41111111110	(	adb41111111110,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m000011_0	),
Adb41111111111	(	adb41111111111,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m000011_0	),
       Adb500(adb500,n0011,n0010,n0009,dbv1),
       Adb501(adb501,n0011,n0010,m0009,m0015),
       Adb510(adb510,n0011,m0010,n0009,dbv1),
       Adb511(adb511,n0011,m0010,m0009,dbv0),
Adb50000000000	(	adb50000000000,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m111010_0	),
Adb50000000001	(	adb50000000001,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m111010_0	),
Adb50000000010	(	adb50000000010,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m111010_0	),
Adb50000000011	(	adb50000000011,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m111010_0	),
Adb50000000100	(	adb50000000100,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m111010_0	),
Adb50000000101	(	adb50000000101,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m111010_0	),
Adb50000000110	(	adb50000000110,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m111010_0	),
Adb50000000111	(	adb50000000111,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m111010_0	),
Adb50000001000	(	adb50000001000,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m111010_0	),
Adb50000001001	(	adb50000001001,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m111010_0	),
Adb50000001010	(	adb50000001010,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m111010_0	),
Adb50000001011	(	adb50000001011,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m111010_0	),
Adb50000001100	(	adb50000001100,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m111010_0	),
Adb50000001101	(	adb50000001101,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m111010_0	),
Adb50000001110	(	adb50000001110,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m111010_0	),
Adb50000001111	(	adb50000001111,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m111010_0	),
Adb50000010000	(	adb50000010000,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m111010_0	),
Adb50000010001	(	adb50000010001,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m111010_0	),
Adb50000010010	(	adb50000010010,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m111010_0	),
Adb50000010011	(	adb50000010011,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m111010_0	),
Adb50000010100	(	adb50000010100,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m111010_0	),
Adb50000010101	(	adb50000010101,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m111010_0	),
Adb50000010110	(	adb50000010110,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m111010_0	),
Adb50000010111	(	adb50000010111,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m111010_0	),
Adb50000011000	(	adb50000011000,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m111010_0	),
Adb50000011001	(	adb50000011001,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m111010_0	),
Adb50000011010	(	adb50000011010,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m111010_0	),
Adb50000011011	(	adb50000011011,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m111010_0	),
Adb50000011100	(	adb50000011100,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m111010_0	),
Adb50000011101	(	adb50000011101,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m111010_0	),
Adb50000011110	(	adb50000011110,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m111010_0	),
Adb50000011111	(	adb50000011111,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m111010_0	),
Adb50000100000	(	adb50000100000,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m111010_0	),
Adb50000100001	(	adb50000100001,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m111010_0	),
Adb50000100010	(	adb50000100010,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m111010_0	),
Adb50000100011	(	adb50000100011,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m111010_0	),
Adb50000100100	(	adb50000100100,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m111010_0	),
Adb50000100101	(	adb50000100101,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m111010_0	),
Adb50000100110	(	adb50000100110,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m111010_0	),
Adb50000100111	(	adb50000100111,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m111010_0	),
Adb50000101000	(	adb50000101000,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m111010_0	),
Adb50000101001	(	adb50000101001,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m111010_0	),
Adb50000101010	(	adb50000101010,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m111010_0	),
Adb50000101011	(	adb50000101011,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m111010_0	),
Adb50000101100	(	adb50000101100,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m111010_0	),
Adb50000101101	(	adb50000101101,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m111010_0	),
Adb50000101110	(	adb50000101110,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m111010_0	),
Adb50000101111	(	adb50000101111,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m111010_0	),
Adb50000110000	(	adb50000110000,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m111010_0	),
Adb50000110001	(	adb50000110001,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m111010_0	),
Adb50000110010	(	adb50000110010,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m111010_0	),
Adb50000110011	(	adb50000110011,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m111010_0	),
Adb50000110100	(	adb50000110100,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m111010_0	),
Adb50000110101	(	adb50000110101,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m111010_0	),
Adb50000110110	(	adb50000110110,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m111010_0	),
Adb50000110111	(	adb50000110111,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m111010_0	),
Adb50000111000	(	adb50000111000,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m111010_0	),
Adb50000111001	(	adb50000111001,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m111010_0	),
Adb50000111010	(	adb50000111010,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m111010_0	),
Adb50000111011	(	adb50000111011,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m111010_0	),
Adb50000111100	(	adb50000111100,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m111010_0	),
Adb50000111101	(	adb50000111101,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m111010_0	),
Adb50000111110	(	adb50000111110,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m111010_0	),
Adb50000111111	(	adb50000111111,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m111010_0	),
Adb50001000000	(	adb50001000000,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m111010_0	),
Adb50001000001	(	adb50001000001,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m111010_0	),
Adb50001000010	(	adb50001000010,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m111010_0	),
Adb50001000011	(	adb50001000011,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m111010_0	),
Adb50001000100	(	adb50001000100,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m111010_0	),
Adb50001000101	(	adb50001000101,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m111010_0	),
Adb50001000110	(	adb50001000110,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m111010_0	),
Adb50001000111	(	adb50001000111,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m111010_0	),
Adb50001001000	(	adb50001001000,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m111010_0	),
Adb50001001001	(	adb50001001001,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m111010_0	),
Adb50001001010	(	adb50001001010,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m111010_0	),
Adb50001001011	(	adb50001001011,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m111010_0	),
Adb50001001100	(	adb50001001100,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m111010_0	),
Adb50001001101	(	adb50001001101,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m111010_0	),
Adb50001001110	(	adb50001001110,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m111010_0	),
Adb50001001111	(	adb50001001111,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m111010_0	),
Adb50001010000	(	adb50001010000,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m111010_0	),
Adb50001010001	(	adb50001010001,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m111010_0	),
Adb50001010010	(	adb50001010010,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m111010_0	),
Adb50001010011	(	adb50001010011,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m111010_0	),
Adb50001010100	(	adb50001010100,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m111010_0	),
Adb50001010101	(	adb50001010101,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m111010_0	),
Adb50001010110	(	adb50001010110,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m111010_0	),
Adb50001010111	(	adb50001010111,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m111010_0	),
Adb50001011000	(	adb50001011000,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m111010_0	),
Adb50001011001	(	adb50001011001,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m111010_0	),
Adb50001011010	(	adb50001011010,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m111010_0	),
Adb50001011011	(	adb50001011011,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m111010_0	),
Adb50001011100	(	adb50001011100,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m111010_0	),
Adb50001011101	(	adb50001011101,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m111010_0	),
Adb50001011110	(	adb50001011110,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m111010_0	),
Adb50001011111	(	adb50001011111,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m111010_0	),
Adb50001100000	(	adb50001100000,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m111010_0	),
Adb50001100001	(	adb50001100001,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m111010_0	),
Adb50001100010	(	adb50001100010,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m111010_0	),
Adb50001100011	(	adb50001100011,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m111010_0	),
Adb50001100100	(	adb50001100100,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m111010_0	),
Adb50001100101	(	adb50001100101,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m111010_0	),
Adb50001100110	(	adb50001100110,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m111010_0	),
Adb50001100111	(	adb50001100111,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m111010_0	),
Adb50001101000	(	adb50001101000,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m111010_0	),
Adb50001101001	(	adb50001101001,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m111010_0	),
Adb50001101010	(	adb50001101010,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m111010_0	),
Adb50001101011	(	adb50001101011,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m111010_0	),
Adb50001101100	(	adb50001101100,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m111010_0	),
Adb50001101101	(	adb50001101101,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m111010_0	),
Adb50001101110	(	adb50001101110,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m111010_0	),
Adb50001101111	(	adb50001101111,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m111010_0	),
Adb50001110000	(	adb50001110000,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m111010_0	),
Adb50001110001	(	adb50001110001,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m111010_0	),
Adb50001110010	(	adb50001110010,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m111010_0	),
Adb50001110011	(	adb50001110011,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m111010_0	),
Adb50001110100	(	adb50001110100,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m111010_0	),
Adb50001110101	(	adb50001110101,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m111010_0	),
Adb50001110110	(	adb50001110110,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m111010_0	),
Adb50001110111	(	adb50001110111,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m111010_0	),
Adb50001111000	(	adb50001111000,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m111010_0	),
Adb50001111001	(	adb50001111001,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m111010_0	),
Adb50001111010	(	adb50001111010,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m111010_0	),
Adb50001111011	(	adb50001111011,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m111010_0	),
Adb50001111100	(	adb50001111100,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m111010_0	),
Adb50001111101	(	adb50001111101,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m111010_0	),
Adb50001111110	(	adb50001111110,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m111010_0	),
Adb50001111111	(	adb50001111111,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m111010_0	),
Adb50010000000	(	adb50010000000,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m110010_0	),
Adb50010000001	(	adb50010000001,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m110010_0	),
Adb50010000010	(	adb50010000010,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m110010_0	),
Adb50010000011	(	adb50010000011,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m110010_0	),
Adb50010000100	(	adb50010000100,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m110010_0	),
Adb50010000101	(	adb50010000101,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m110010_0	),
Adb50010000110	(	adb50010000110,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m110010_0	),
Adb50010000111	(	adb50010000111,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m110010_0	),
Adb50010001000	(	adb50010001000,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m110010_0	),
Adb50010001001	(	adb50010001001,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m110010_0	),
Adb50010001010	(	adb50010001010,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m110010_0	),
Adb50010001011	(	adb50010001011,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m110010_0	),
Adb50010001100	(	adb50010001100,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m110010_0	),
Adb50010001101	(	adb50010001101,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m110010_0	),
Adb50010001110	(	adb50010001110,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m110010_0	),
Adb50010001111	(	adb50010001111,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m110010_0	),
Adb50010010000	(	adb50010010000,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m110010_0	),
Adb50010010001	(	adb50010010001,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m110010_0	),
Adb50010010010	(	adb50010010010,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m110010_0	),
Adb50010010011	(	adb50010010011,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m110010_0	),
Adb50010010100	(	adb50010010100,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m110010_0	),
Adb50010010101	(	adb50010010101,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m110010_0	),
Adb50010010110	(	adb50010010110,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m110010_0	),
Adb50010010111	(	adb50010010111,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m110010_0	),
Adb50010011000	(	adb50010011000,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m110010_0	),
Adb50010011001	(	adb50010011001,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m110010_0	),
Adb50010011010	(	adb50010011010,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m110010_0	),
Adb50010011011	(	adb50010011011,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m110010_0	),
Adb50010011100	(	adb50010011100,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m110010_0	),
Adb50010011101	(	adb50010011101,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m110010_0	),
Adb50010011110	(	adb50010011110,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m110010_0	),
Adb50010011111	(	adb50010011111,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m110010_0	),
Adb50010100000	(	adb50010100000,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m110010_0	),
Adb50010100001	(	adb50010100001,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m110010_0	),
Adb50010100010	(	adb50010100010,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m110010_0	),
Adb50010100011	(	adb50010100011,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m110010_0	),
Adb50010100100	(	adb50010100100,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m110010_0	),
Adb50010100101	(	adb50010100101,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m110010_0	),
Adb50010100110	(	adb50010100110,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m110010_0	),
Adb50010100111	(	adb50010100111,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m110010_0	),
Adb50010101000	(	adb50010101000,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m110010_0	),
Adb50010101001	(	adb50010101001,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m110010_0	),
Adb50010101010	(	adb50010101010,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m110010_0	),
Adb50010101011	(	adb50010101011,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m110010_0	),
Adb50010101100	(	adb50010101100,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m110010_0	),
Adb50010101101	(	adb50010101101,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m110010_0	),
Adb50010101110	(	adb50010101110,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m110010_0	),
Adb50010101111	(	adb50010101111,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m110010_0	),
Adb50010110000	(	adb50010110000,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m110010_0	),
Adb50010110001	(	adb50010110001,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m110010_0	),
Adb50010110010	(	adb50010110010,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m110010_0	),
Adb50010110011	(	adb50010110011,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m110010_0	),
Adb50010110100	(	adb50010110100,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m110010_0	),
Adb50010110101	(	adb50010110101,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m110010_0	),
Adb50010110110	(	adb50010110110,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m110010_0	),
Adb50010110111	(	adb50010110111,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m110010_0	),
Adb50010111000	(	adb50010111000,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m110010_0	),
Adb50010111001	(	adb50010111001,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m110010_0	),
Adb50010111010	(	adb50010111010,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m110010_0	),
Adb50010111011	(	adb50010111011,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m110010_0	),
Adb50010111100	(	adb50010111100,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m110010_0	),
Adb50010111101	(	adb50010111101,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m110010_0	),
Adb50010111110	(	adb50010111110,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m110010_0	),
Adb50010111111	(	adb50010111111,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m110010_0	),
Adb50011000000	(	adb50011000000,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m110010_0	),
Adb50011000001	(	adb50011000001,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m110010_0	),
Adb50011000010	(	adb50011000010,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m110010_0	),
Adb50011000011	(	adb50011000011,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m110010_0	),
Adb50011000100	(	adb50011000100,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m110010_0	),
Adb50011000101	(	adb50011000101,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m110010_0	),
Adb50011000110	(	adb50011000110,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m110010_0	),
Adb50011000111	(	adb50011000111,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m110010_0	),
Adb50011001000	(	adb50011001000,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m110010_0	),
Adb50011001001	(	adb50011001001,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m110010_0	),
Adb50011001010	(	adb50011001010,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m110010_0	),
Adb50011001011	(	adb50011001011,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m110010_0	),
Adb50011001100	(	adb50011001100,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m110010_0	),
Adb50011001101	(	adb50011001101,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m110010_0	),
Adb50011001110	(	adb50011001110,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m110010_0	),
Adb50011001111	(	adb50011001111,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m110010_0	),
Adb50011010000	(	adb50011010000,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m110010_0	),
Adb50011010001	(	adb50011010001,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m110010_0	),
Adb50011010010	(	adb50011010010,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m110010_0	),
Adb50011010011	(	adb50011010011,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m110010_0	),
Adb50011010100	(	adb50011010100,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m110010_0	),
Adb50011010101	(	adb50011010101,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m110010_0	),
Adb50011010110	(	adb50011010110,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m110010_0	),
Adb50011010111	(	adb50011010111,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m110010_0	),
Adb50011011000	(	adb50011011000,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m110010_0	),
Adb50011011001	(	adb50011011001,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m110010_0	),
Adb50011011010	(	adb50011011010,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m110010_0	),
Adb50011011011	(	adb50011011011,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m110010_0	),
Adb50011011100	(	adb50011011100,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m110010_0	),
Adb50011011101	(	adb50011011101,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m110010_0	),
Adb50011011110	(	adb50011011110,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m110010_0	),
Adb50011011111	(	adb50011011111,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m110010_0	),
Adb50011100000	(	adb50011100000,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m110010_0	),
Adb50011100001	(	adb50011100001,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m110010_0	),
Adb50011100010	(	adb50011100010,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m110010_0	),
Adb50011100011	(	adb50011100011,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m110010_0	),
Adb50011100100	(	adb50011100100,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m110010_0	),
Adb50011100101	(	adb50011100101,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m110010_0	),
Adb50011100110	(	adb50011100110,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m110010_0	),
Adb50011100111	(	adb50011100111,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m110010_0	),
Adb50011101000	(	adb50011101000,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m110010_0	),
Adb50011101001	(	adb50011101001,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m110010_0	),
Adb50011101010	(	adb50011101010,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m110010_0	),
Adb50011101011	(	adb50011101011,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m110010_0	),
Adb50011101100	(	adb50011101100,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m110010_0	),
Adb50011101101	(	adb50011101101,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m110010_0	),
Adb50011101110	(	adb50011101110,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m110010_0	),
Adb50011101111	(	adb50011101111,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m110010_0	),
Adb50011110000	(	adb50011110000,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m110010_0	),
Adb50011110001	(	adb50011110001,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m110010_0	),
Adb50011110010	(	adb50011110010,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m110010_0	),
Adb50011110011	(	adb50011110011,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m110010_0	),
Adb50011110100	(	adb50011110100,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m110010_0	),
Adb50011110101	(	adb50011110101,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m110010_0	),
Adb50011110110	(	adb50011110110,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m110010_0	),
Adb50011110111	(	adb50011110111,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m110010_0	),
Adb50011111000	(	adb50011111000,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m110010_0	),
Adb50011111001	(	adb50011111001,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m110010_0	),
Adb50011111010	(	adb50011111010,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m110010_0	),
Adb50011111011	(	adb50011111011,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m110010_0	),
Adb50011111100	(	adb50011111100,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m110010_0	),
Adb50011111101	(	adb50011111101,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m110010_0	),
Adb50011111110	(	adb50011111110,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m110010_0	),
Adb50011111111	(	adb50011111111,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m110010_0	),
Adb50100000000	(	adb50100000000,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m101010_0	),
Adb50100000001	(	adb50100000001,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m101010_0	),
Adb50100000010	(	adb50100000010,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m101010_0	),
Adb50100000011	(	adb50100000011,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m101010_0	),
Adb50100000100	(	adb50100000100,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m101010_0	),
Adb50100000101	(	adb50100000101,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m101010_0	),
Adb50100000110	(	adb50100000110,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m101010_0	),
Adb50100000111	(	adb50100000111,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m101010_0	),
Adb50100001000	(	adb50100001000,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m101010_0	),
Adb50100001001	(	adb50100001001,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m101010_0	),
Adb50100001010	(	adb50100001010,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m101010_0	),
Adb50100001011	(	adb50100001011,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m101010_0	),
Adb50100001100	(	adb50100001100,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m101010_0	),
Adb50100001101	(	adb50100001101,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m101010_0	),
Adb50100001110	(	adb50100001110,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m101010_0	),
Adb50100001111	(	adb50100001111,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m101010_0	),
Adb50100010000	(	adb50100010000,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m101010_0	),
Adb50100010001	(	adb50100010001,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m101010_0	),
Adb50100010010	(	adb50100010010,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m101010_0	),
Adb50100010011	(	adb50100010011,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m101010_0	),
Adb50100010100	(	adb50100010100,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m101010_0	),
Adb50100010101	(	adb50100010101,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m101010_0	),
Adb50100010110	(	adb50100010110,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m101010_0	),
Adb50100010111	(	adb50100010111,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m101010_0	),
Adb50100011000	(	adb50100011000,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m101010_0	),
Adb50100011001	(	adb50100011001,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m101010_0	),
Adb50100011010	(	adb50100011010,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m101010_0	),
Adb50100011011	(	adb50100011011,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m101010_0	),
Adb50100011100	(	adb50100011100,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m101010_0	),
Adb50100011101	(	adb50100011101,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m101010_0	),
Adb50100011110	(	adb50100011110,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m101010_0	),
Adb50100011111	(	adb50100011111,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m101010_0	),
Adb50100100000	(	adb50100100000,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m101010_0	),
Adb50100100001	(	adb50100100001,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m101010_0	),
Adb50100100010	(	adb50100100010,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m101010_0	),
Adb50100100011	(	adb50100100011,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m101010_0	),
Adb50100100100	(	adb50100100100,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m101010_0	),
Adb50100100101	(	adb50100100101,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m101010_0	),
Adb50100100110	(	adb50100100110,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m101010_0	),
Adb50100100111	(	adb50100100111,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m101010_0	),
Adb50100101000	(	adb50100101000,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m101010_0	),
Adb50100101001	(	adb50100101001,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m101010_0	),
Adb50100101010	(	adb50100101010,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m101010_0	),
Adb50100101011	(	adb50100101011,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m101010_0	),
Adb50100101100	(	adb50100101100,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m101010_0	),
Adb50100101101	(	adb50100101101,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m101010_0	),
Adb50100101110	(	adb50100101110,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m101010_0	),
Adb50100101111	(	adb50100101111,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m101010_0	),
Adb50100110000	(	adb50100110000,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m101010_0	),
Adb50100110001	(	adb50100110001,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m101010_0	),
Adb50100110010	(	adb50100110010,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m101010_0	),
Adb50100110011	(	adb50100110011,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m101010_0	),
Adb50100110100	(	adb50100110100,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m101010_0	),
Adb50100110101	(	adb50100110101,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m101010_0	),
Adb50100110110	(	adb50100110110,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m101010_0	),
Adb50100110111	(	adb50100110111,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m101010_0	),
Adb50100111000	(	adb50100111000,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m101010_0	),
Adb50100111001	(	adb50100111001,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m101010_0	),
Adb50100111010	(	adb50100111010,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m101010_0	),
Adb50100111011	(	adb50100111011,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m101010_0	),
Adb50100111100	(	adb50100111100,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m101010_0	),
Adb50100111101	(	adb50100111101,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m101010_0	),
Adb50100111110	(	adb50100111110,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m101010_0	),
Adb50100111111	(	adb50100111111,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m101010_0	),
Adb50101000000	(	adb50101000000,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m101010_0	),
Adb50101000001	(	adb50101000001,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m101010_0	),
Adb50101000010	(	adb50101000010,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m101010_0	),
Adb50101000011	(	adb50101000011,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m101010_0	),
Adb50101000100	(	adb50101000100,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m101010_0	),
Adb50101000101	(	adb50101000101,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m101010_0	),
Adb50101000110	(	adb50101000110,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m101010_0	),
Adb50101000111	(	adb50101000111,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m101010_0	),
Adb50101001000	(	adb50101001000,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m101010_0	),
Adb50101001001	(	adb50101001001,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m101010_0	),
Adb50101001010	(	adb50101001010,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m101010_0	),
Adb50101001011	(	adb50101001011,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m101010_0	),
Adb50101001100	(	adb50101001100,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m101010_0	),
Adb50101001101	(	adb50101001101,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m101010_0	),
Adb50101001110	(	adb50101001110,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m101010_0	),
Adb50101001111	(	adb50101001111,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m101010_0	),
Adb50101010000	(	adb50101010000,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m101010_0	),
Adb50101010001	(	adb50101010001,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m101010_0	),
Adb50101010010	(	adb50101010010,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m101010_0	),
Adb50101010011	(	adb50101010011,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m101010_0	),
Adb50101010100	(	adb50101010100,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m101010_0	),
Adb50101010101	(	adb50101010101,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m101010_0	),
Adb50101010110	(	adb50101010110,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m101010_0	),
Adb50101010111	(	adb50101010111,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m101010_0	),
Adb50101011000	(	adb50101011000,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m101010_0	),
Adb50101011001	(	adb50101011001,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m101010_0	),
Adb50101011010	(	adb50101011010,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m101010_0	),
Adb50101011011	(	adb50101011011,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m101010_0	),
Adb50101011100	(	adb50101011100,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m101010_0	),
Adb50101011101	(	adb50101011101,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m101010_0	),
Adb50101011110	(	adb50101011110,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m101010_0	),
Adb50101011111	(	adb50101011111,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m101010_0	),
Adb50101100000	(	adb50101100000,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m101010_0	),
Adb50101100001	(	adb50101100001,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m101010_0	),
Adb50101100010	(	adb50101100010,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m101010_0	),
Adb50101100011	(	adb50101100011,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m101010_0	),
Adb50101100100	(	adb50101100100,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m101010_0	),
Adb50101100101	(	adb50101100101,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m101010_0	),
Adb50101100110	(	adb50101100110,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m101010_0	),
Adb50101100111	(	adb50101100111,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m101010_0	),
Adb50101101000	(	adb50101101000,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m101010_0	),
Adb50101101001	(	adb50101101001,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m101010_0	),
Adb50101101010	(	adb50101101010,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m101010_0	),
Adb50101101011	(	adb50101101011,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m101010_0	),
Adb50101101100	(	adb50101101100,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m101010_0	),
Adb50101101101	(	adb50101101101,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m101010_0	),
Adb50101101110	(	adb50101101110,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m101010_0	),
Adb50101101111	(	adb50101101111,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m101010_0	),
Adb50101110000	(	adb50101110000,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m101010_0	),
Adb50101110001	(	adb50101110001,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m101010_0	),
Adb50101110010	(	adb50101110010,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m101010_0	),
Adb50101110011	(	adb50101110011,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m101010_0	),
Adb50101110100	(	adb50101110100,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m101010_0	),
Adb50101110101	(	adb50101110101,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m101010_0	),
Adb50101110110	(	adb50101110110,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m101010_0	),
Adb50101110111	(	adb50101110111,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m101010_0	),
Adb50101111000	(	adb50101111000,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m101010_0	),
Adb50101111001	(	adb50101111001,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m101010_0	),
Adb50101111010	(	adb50101111010,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m101010_0	),
Adb50101111011	(	adb50101111011,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m101010_0	),
Adb50101111100	(	adb50101111100,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m101010_0	),
Adb50101111101	(	adb50101111101,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m101010_0	),
Adb50101111110	(	adb50101111110,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m101010_0	),
Adb50101111111	(	adb50101111111,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m101010_0	),
Adb50110000000	(	adb50110000000,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m100010_0	),
Adb50110000001	(	adb50110000001,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m100010_0	),
Adb50110000010	(	adb50110000010,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m100010_0	),
Adb50110000011	(	adb50110000011,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m100010_0	),
Adb50110000100	(	adb50110000100,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m100010_0	),
Adb50110000101	(	adb50110000101,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m100010_0	),
Adb50110000110	(	adb50110000110,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m100010_0	),
Adb50110000111	(	adb50110000111,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m100010_0	),
Adb50110001000	(	adb50110001000,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m100010_0	),
Adb50110001001	(	adb50110001001,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m100010_0	),
Adb50110001010	(	adb50110001010,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m100010_0	),
Adb50110001011	(	adb50110001011,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m100010_0	),
Adb50110001100	(	adb50110001100,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m100010_0	),
Adb50110001101	(	adb50110001101,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m100010_0	),
Adb50110001110	(	adb50110001110,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m100010_0	),
Adb50110001111	(	adb50110001111,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m100010_0	),
Adb50110010000	(	adb50110010000,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m100010_0	),
Adb50110010001	(	adb50110010001,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m100010_0	),
Adb50110010010	(	adb50110010010,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m100010_0	),
Adb50110010011	(	adb50110010011,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m100010_0	),
Adb50110010100	(	adb50110010100,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m100010_0	),
Adb50110010101	(	adb50110010101,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m100010_0	),
Adb50110010110	(	adb50110010110,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m100010_0	),
Adb50110010111	(	adb50110010111,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m100010_0	),
Adb50110011000	(	adb50110011000,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m100010_0	),
Adb50110011001	(	adb50110011001,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m100010_0	),
Adb50110011010	(	adb50110011010,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m100010_0	),
Adb50110011011	(	adb50110011011,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m100010_0	),
Adb50110011100	(	adb50110011100,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m100010_0	),
Adb50110011101	(	adb50110011101,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m100010_0	),
Adb50110011110	(	adb50110011110,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m100010_0	),
Adb50110011111	(	adb50110011111,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m100010_0	),
Adb50110100000	(	adb50110100000,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m100010_0	),
Adb50110100001	(	adb50110100001,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m100010_0	),
Adb50110100010	(	adb50110100010,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m100010_0	),
Adb50110100011	(	adb50110100011,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m100010_0	),
Adb50110100100	(	adb50110100100,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m100010_0	),
Adb50110100101	(	adb50110100101,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m100010_0	),
Adb50110100110	(	adb50110100110,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m100010_0	),
Adb50110100111	(	adb50110100111,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m100010_0	),
Adb50110101000	(	adb50110101000,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m100010_0	),
Adb50110101001	(	adb50110101001,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m100010_0	),
Adb50110101010	(	adb50110101010,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m100010_0	),
Adb50110101011	(	adb50110101011,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m100010_0	),
Adb50110101100	(	adb50110101100,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m100010_0	),
Adb50110101101	(	adb50110101101,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m100010_0	),
Adb50110101110	(	adb50110101110,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m100010_0	),
Adb50110101111	(	adb50110101111,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m100010_0	),
Adb50110110000	(	adb50110110000,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m100010_0	),
Adb50110110001	(	adb50110110001,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m100010_0	),
Adb50110110010	(	adb50110110010,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m100010_0	),
Adb50110110011	(	adb50110110011,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m100010_0	),
Adb50110110100	(	adb50110110100,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m100010_0	),
Adb50110110101	(	adb50110110101,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m100010_0	),
Adb50110110110	(	adb50110110110,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m100010_0	),
Adb50110110111	(	adb50110110111,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m100010_0	),
Adb50110111000	(	adb50110111000,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m100010_0	),
Adb50110111001	(	adb50110111001,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m100010_0	),
Adb50110111010	(	adb50110111010,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m100010_0	),
Adb50110111011	(	adb50110111011,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m100010_0	),
Adb50110111100	(	adb50110111100,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m100010_0	),
Adb50110111101	(	adb50110111101,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m100010_0	),
Adb50110111110	(	adb50110111110,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m100010_0	),
Adb50110111111	(	adb50110111111,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m100010_0	),
Adb50111000000	(	adb50111000000,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m100010_0	),
Adb50111000001	(	adb50111000001,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m100010_0	),
Adb50111000010	(	adb50111000010,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m100010_0	),
Adb50111000011	(	adb50111000011,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m100010_0	),
Adb50111000100	(	adb50111000100,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m100010_0	),
Adb50111000101	(	adb50111000101,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m100010_0	),
Adb50111000110	(	adb50111000110,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m100010_0	),
Adb50111000111	(	adb50111000111,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m100010_0	),
Adb50111001000	(	adb50111001000,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m100010_0	),
Adb50111001001	(	adb50111001001,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m100010_0	),
Adb50111001010	(	adb50111001010,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m100010_0	),
Adb50111001011	(	adb50111001011,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m100010_0	),
Adb50111001100	(	adb50111001100,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m100010_0	),
Adb50111001101	(	adb50111001101,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m100010_0	),
Adb50111001110	(	adb50111001110,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m100010_0	),
Adb50111001111	(	adb50111001111,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m100010_0	),
Adb50111010000	(	adb50111010000,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m100010_0	),
Adb50111010001	(	adb50111010001,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m100010_0	),
Adb50111010010	(	adb50111010010,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m100010_0	),
Adb50111010011	(	adb50111010011,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m100010_0	),
Adb50111010100	(	adb50111010100,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m100010_0	),
Adb50111010101	(	adb50111010101,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m100010_0	),
Adb50111010110	(	adb50111010110,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m100010_0	),
Adb50111010111	(	adb50111010111,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m100010_0	),
Adb50111011000	(	adb50111011000,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m100010_0	),
Adb50111011001	(	adb50111011001,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m100010_0	),
Adb50111011010	(	adb50111011010,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m100010_0	),
Adb50111011011	(	adb50111011011,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m100010_0	),
Adb50111011100	(	adb50111011100,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m100010_0	),
Adb50111011101	(	adb50111011101,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m100010_0	),
Adb50111011110	(	adb50111011110,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m100010_0	),
Adb50111011111	(	adb50111011111,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m100010_0	),
Adb50111100000	(	adb50111100000,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m100010_0	),
Adb50111100001	(	adb50111100001,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m100010_0	),
Adb50111100010	(	adb50111100010,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m100010_0	),
Adb50111100011	(	adb50111100011,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m100010_0	),
Adb50111100100	(	adb50111100100,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m100010_0	),
Adb50111100101	(	adb50111100101,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m100010_0	),
Adb50111100110	(	adb50111100110,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m100010_0	),
Adb50111100111	(	adb50111100111,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m100010_0	),
Adb50111101000	(	adb50111101000,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m100010_0	),
Adb50111101001	(	adb50111101001,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m100010_0	),
Adb50111101010	(	adb50111101010,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m100010_0	),
Adb50111101011	(	adb50111101011,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m100010_0	),
Adb50111101100	(	adb50111101100,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m100010_0	),
Adb50111101101	(	adb50111101101,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m100010_0	),
Adb50111101110	(	adb50111101110,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m100010_0	),
Adb50111101111	(	adb50111101111,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m100010_0	),
Adb50111110000	(	adb50111110000,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m100010_0	),
Adb50111110001	(	adb50111110001,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m100010_0	),
Adb50111110010	(	adb50111110010,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m100010_0	),
Adb50111110011	(	adb50111110011,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m100010_0	),
Adb50111110100	(	adb50111110100,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m100010_0	),
Adb50111110101	(	adb50111110101,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m100010_0	),
Adb50111110110	(	adb50111110110,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m100010_0	),
Adb50111110111	(	adb50111110111,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m100010_0	),
Adb50111111000	(	adb50111111000,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m100010_0	),
Adb50111111001	(	adb50111111001,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m100010_0	),
Adb50111111010	(	adb50111111010,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m100010_0	),
Adb50111111011	(	adb50111111011,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m100010_0	),
Adb50111111100	(	adb50111111100,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m100010_0	),
Adb50111111101	(	adb50111111101,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m100010_0	),
Adb50111111110	(	adb50111111110,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m100010_0	),
Adb50111111111	(	adb50111111111,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m100010_0	),
Adb51000000000	(	adb51000000000,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m011010_0	),
Adb51000000001	(	adb51000000001,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m011010_0	),
Adb51000000010	(	adb51000000010,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m011010_0	),
Adb51000000011	(	adb51000000011,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m011010_0	),
Adb51000000100	(	adb51000000100,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m011010_0	),
Adb51000000101	(	adb51000000101,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m011010_0	),
Adb51000000110	(	adb51000000110,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m011010_0	),
Adb51000000111	(	adb51000000111,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m011010_0	),
Adb51000001000	(	adb51000001000,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m011010_0	),
Adb51000001001	(	adb51000001001,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m011010_0	),
Adb51000001010	(	adb51000001010,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m011010_0	),
Adb51000001011	(	adb51000001011,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m011010_0	),
Adb51000001100	(	adb51000001100,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m011010_0	),
Adb51000001101	(	adb51000001101,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m011010_0	),
Adb51000001110	(	adb51000001110,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m011010_0	),
Adb51000001111	(	adb51000001111,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m011010_0	),
Adb51000010000	(	adb51000010000,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m011010_0	),
Adb51000010001	(	adb51000010001,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m011010_0	),
Adb51000010010	(	adb51000010010,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m011010_0	),
Adb51000010011	(	adb51000010011,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m011010_0	),
Adb51000010100	(	adb51000010100,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m011010_0	),
Adb51000010101	(	adb51000010101,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m011010_0	),
Adb51000010110	(	adb51000010110,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m011010_0	),
Adb51000010111	(	adb51000010111,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m011010_0	),
Adb51000011000	(	adb51000011000,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m011010_0	),
Adb51000011001	(	adb51000011001,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m011010_0	),
Adb51000011010	(	adb51000011010,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m011010_0	),
Adb51000011011	(	adb51000011011,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m011010_0	),
Adb51000011100	(	adb51000011100,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m011010_0	),
Adb51000011101	(	adb51000011101,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m011010_0	),
Adb51000011110	(	adb51000011110,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m011010_0	),
Adb51000011111	(	adb51000011111,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m011010_0	),
Adb51000100000	(	adb51000100000,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m011010_0	),
Adb51000100001	(	adb51000100001,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m011010_0	),
Adb51000100010	(	adb51000100010,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m011010_0	),
Adb51000100011	(	adb51000100011,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m011010_0	),
Adb51000100100	(	adb51000100100,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m011010_0	),
Adb51000100101	(	adb51000100101,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m011010_0	),
Adb51000100110	(	adb51000100110,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m011010_0	),
Adb51000100111	(	adb51000100111,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m011010_0	),
Adb51000101000	(	adb51000101000,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m011010_0	),
Adb51000101001	(	adb51000101001,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m011010_0	),
Adb51000101010	(	adb51000101010,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m011010_0	),
Adb51000101011	(	adb51000101011,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m011010_0	),
Adb51000101100	(	adb51000101100,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m011010_0	),
Adb51000101101	(	adb51000101101,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m011010_0	),
Adb51000101110	(	adb51000101110,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m011010_0	),
Adb51000101111	(	adb51000101111,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m011010_0	),
Adb51000110000	(	adb51000110000,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m011010_0	),
Adb51000110001	(	adb51000110001,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m011010_0	),
Adb51000110010	(	adb51000110010,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m011010_0	),
Adb51000110011	(	adb51000110011,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m011010_0	),
Adb51000110100	(	adb51000110100,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m011010_0	),
Adb51000110101	(	adb51000110101,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m011010_0	),
Adb51000110110	(	adb51000110110,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m011010_0	),
Adb51000110111	(	adb51000110111,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m011010_0	),
Adb51000111000	(	adb51000111000,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m011010_0	),
Adb51000111001	(	adb51000111001,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m011010_0	),
Adb51000111010	(	adb51000111010,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m011010_0	),
Adb51000111011	(	adb51000111011,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m011010_0	),
Adb51000111100	(	adb51000111100,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m011010_0	),
Adb51000111101	(	adb51000111101,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m011010_0	),
Adb51000111110	(	adb51000111110,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m011010_0	),
Adb51000111111	(	adb51000111111,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m011010_0	),
Adb51001000000	(	adb51001000000,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m011010_0	),
Adb51001000001	(	adb51001000001,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m011010_0	),
Adb51001000010	(	adb51001000010,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m011010_0	),
Adb51001000011	(	adb51001000011,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m011010_0	),
Adb51001000100	(	adb51001000100,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m011010_0	),
Adb51001000101	(	adb51001000101,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m011010_0	),
Adb51001000110	(	adb51001000110,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m011010_0	),
Adb51001000111	(	adb51001000111,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m011010_0	),
Adb51001001000	(	adb51001001000,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m011010_0	),
Adb51001001001	(	adb51001001001,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m011010_0	),
Adb51001001010	(	adb51001001010,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m011010_0	),
Adb51001001011	(	adb51001001011,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m011010_0	),
Adb51001001100	(	adb51001001100,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m011010_0	),
Adb51001001101	(	adb51001001101,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m011010_0	),
Adb51001001110	(	adb51001001110,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m011010_0	),
Adb51001001111	(	adb51001001111,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m011010_0	),
Adb51001010000	(	adb51001010000,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m011010_0	),
Adb51001010001	(	adb51001010001,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m011010_0	),
Adb51001010010	(	adb51001010010,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m011010_0	),
Adb51001010011	(	adb51001010011,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m011010_0	),
Adb51001010100	(	adb51001010100,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m011010_0	),
Adb51001010101	(	adb51001010101,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m011010_0	),
Adb51001010110	(	adb51001010110,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m011010_0	),
Adb51001010111	(	adb51001010111,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m011010_0	),
Adb51001011000	(	adb51001011000,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m011010_0	),
Adb51001011001	(	adb51001011001,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m011010_0	),
Adb51001011010	(	adb51001011010,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m011010_0	),
Adb51001011011	(	adb51001011011,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m011010_0	),
Adb51001011100	(	adb51001011100,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m011010_0	),
Adb51001011101	(	adb51001011101,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m011010_0	),
Adb51001011110	(	adb51001011110,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m011010_0	),
Adb51001011111	(	adb51001011111,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m011010_0	),
Adb51001100000	(	adb51001100000,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m011010_0	),
Adb51001100001	(	adb51001100001,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m011010_0	),
Adb51001100010	(	adb51001100010,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m011010_0	),
Adb51001100011	(	adb51001100011,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m011010_0	),
Adb51001100100	(	adb51001100100,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m011010_0	),
Adb51001100101	(	adb51001100101,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m011010_0	),
Adb51001100110	(	adb51001100110,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m011010_0	),
Adb51001100111	(	adb51001100111,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m011010_0	),
Adb51001101000	(	adb51001101000,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m011010_0	),
Adb51001101001	(	adb51001101001,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m011010_0	),
Adb51001101010	(	adb51001101010,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m011010_0	),
Adb51001101011	(	adb51001101011,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m011010_0	),
Adb51001101100	(	adb51001101100,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m011010_0	),
Adb51001101101	(	adb51001101101,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m011010_0	),
Adb51001101110	(	adb51001101110,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m011010_0	),
Adb51001101111	(	adb51001101111,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m011010_0	),
Adb51001110000	(	adb51001110000,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m011010_0	),
Adb51001110001	(	adb51001110001,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m011010_0	),
Adb51001110010	(	adb51001110010,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m011010_0	),
Adb51001110011	(	adb51001110011,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m011010_0	),
Adb51001110100	(	adb51001110100,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m011010_0	),
Adb51001110101	(	adb51001110101,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m011010_0	),
Adb51001110110	(	adb51001110110,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m011010_0	),
Adb51001110111	(	adb51001110111,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m011010_0	),
Adb51001111000	(	adb51001111000,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m011010_0	),
Adb51001111001	(	adb51001111001,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m011010_0	),
Adb51001111010	(	adb51001111010,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m011010_0	),
Adb51001111011	(	adb51001111011,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m011010_0	),
Adb51001111100	(	adb51001111100,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m011010_0	),
Adb51001111101	(	adb51001111101,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m011010_0	),
Adb51001111110	(	adb51001111110,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m011010_0	),
Adb51001111111	(	adb51001111111,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m011010_0	),
Adb51010000000	(	adb51010000000,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m010010_0	),
Adb51010000001	(	adb51010000001,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m010010_0	),
Adb51010000010	(	adb51010000010,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m010010_0	),
Adb51010000011	(	adb51010000011,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m010010_0	),
Adb51010000100	(	adb51010000100,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m010010_0	),
Adb51010000101	(	adb51010000101,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m010010_0	),
Adb51010000110	(	adb51010000110,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m010010_0	),
Adb51010000111	(	adb51010000111,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m010010_0	),
Adb51010001000	(	adb51010001000,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m010010_0	),
Adb51010001001	(	adb51010001001,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m010010_0	),
Adb51010001010	(	adb51010001010,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m010010_0	),
Adb51010001011	(	adb51010001011,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m010010_0	),
Adb51010001100	(	adb51010001100,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m010010_0	),
Adb51010001101	(	adb51010001101,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m010010_0	),
Adb51010001110	(	adb51010001110,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m010010_0	),
Adb51010001111	(	adb51010001111,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m010010_0	),
Adb51010010000	(	adb51010010000,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m010010_0	),
Adb51010010001	(	adb51010010001,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m010010_0	),
Adb51010010010	(	adb51010010010,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m010010_0	),
Adb51010010011	(	adb51010010011,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m010010_0	),
Adb51010010100	(	adb51010010100,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m010010_0	),
Adb51010010101	(	adb51010010101,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m010010_0	),
Adb51010010110	(	adb51010010110,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m010010_0	),
Adb51010010111	(	adb51010010111,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m010010_0	),
Adb51010011000	(	adb51010011000,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m010010_0	),
Adb51010011001	(	adb51010011001,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m010010_0	),
Adb51010011010	(	adb51010011010,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m010010_0	),
Adb51010011011	(	adb51010011011,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m010010_0	),
Adb51010011100	(	adb51010011100,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m010010_0	),
Adb51010011101	(	adb51010011101,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m010010_0	),
Adb51010011110	(	adb51010011110,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m010010_0	),
Adb51010011111	(	adb51010011111,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m010010_0	),
Adb51010100000	(	adb51010100000,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m010010_0	),
Adb51010100001	(	adb51010100001,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m010010_0	),
Adb51010100010	(	adb51010100010,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m010010_0	),
Adb51010100011	(	adb51010100011,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m010010_0	),
Adb51010100100	(	adb51010100100,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m010010_0	),
Adb51010100101	(	adb51010100101,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m010010_0	),
Adb51010100110	(	adb51010100110,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m010010_0	),
Adb51010100111	(	adb51010100111,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m010010_0	),
Adb51010101000	(	adb51010101000,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m010010_0	),
Adb51010101001	(	adb51010101001,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m010010_0	),
Adb51010101010	(	adb51010101010,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m010010_0	),
Adb51010101011	(	adb51010101011,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m010010_0	),
Adb51010101100	(	adb51010101100,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m010010_0	),
Adb51010101101	(	adb51010101101,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m010010_0	),
Adb51010101110	(	adb51010101110,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m010010_0	),
Adb51010101111	(	adb51010101111,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m010010_0	),
Adb51010110000	(	adb51010110000,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m010010_0	),
Adb51010110001	(	adb51010110001,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m010010_0	),
Adb51010110010	(	adb51010110010,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m010010_0	),
Adb51010110011	(	adb51010110011,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m010010_0	),
Adb51010110100	(	adb51010110100,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m010010_0	),
Adb51010110101	(	adb51010110101,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m010010_0	),
Adb51010110110	(	adb51010110110,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m010010_0	),
Adb51010110111	(	adb51010110111,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m010010_0	),
Adb51010111000	(	adb51010111000,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m010010_0	),
Adb51010111001	(	adb51010111001,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m010010_0	),
Adb51010111010	(	adb51010111010,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m010010_0	),
Adb51010111011	(	adb51010111011,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m010010_0	),
Adb51010111100	(	adb51010111100,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m010010_0	),
Adb51010111101	(	adb51010111101,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m010010_0	),
Adb51010111110	(	adb51010111110,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m010010_0	),
Adb51010111111	(	adb51010111111,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m010010_0	),
Adb51011000000	(	adb51011000000,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m010010_0	),
Adb51011000001	(	adb51011000001,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m010010_0	),
Adb51011000010	(	adb51011000010,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m010010_0	),
Adb51011000011	(	adb51011000011,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m010010_0	),
Adb51011000100	(	adb51011000100,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m010010_0	),
Adb51011000101	(	adb51011000101,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m010010_0	),
Adb51011000110	(	adb51011000110,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m010010_0	),
Adb51011000111	(	adb51011000111,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m010010_0	),
Adb51011001000	(	adb51011001000,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m010010_0	),
Adb51011001001	(	adb51011001001,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m010010_0	),
Adb51011001010	(	adb51011001010,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m010010_0	),
Adb51011001011	(	adb51011001011,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m010010_0	),
Adb51011001100	(	adb51011001100,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m010010_0	),
Adb51011001101	(	adb51011001101,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m010010_0	),
Adb51011001110	(	adb51011001110,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m010010_0	),
Adb51011001111	(	adb51011001111,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m010010_0	),
Adb51011010000	(	adb51011010000,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m010010_0	),
Adb51011010001	(	adb51011010001,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m010010_0	),
Adb51011010010	(	adb51011010010,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m010010_0	),
Adb51011010011	(	adb51011010011,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m010010_0	),
Adb51011010100	(	adb51011010100,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m010010_0	),
Adb51011010101	(	adb51011010101,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m010010_0	),
Adb51011010110	(	adb51011010110,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m010010_0	),
Adb51011010111	(	adb51011010111,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m010010_0	),
Adb51011011000	(	adb51011011000,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m010010_0	),
Adb51011011001	(	adb51011011001,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m010010_0	),
Adb51011011010	(	adb51011011010,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m010010_0	),
Adb51011011011	(	adb51011011011,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m010010_0	),
Adb51011011100	(	adb51011011100,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m010010_0	),
Adb51011011101	(	adb51011011101,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m010010_0	),
Adb51011011110	(	adb51011011110,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m010010_0	),
Adb51011011111	(	adb51011011111,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m010010_0	),
Adb51011100000	(	adb51011100000,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m010010_0	),
Adb51011100001	(	adb51011100001,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m010010_0	),
Adb51011100010	(	adb51011100010,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m010010_0	),
Adb51011100011	(	adb51011100011,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m010010_0	),
Adb51011100100	(	adb51011100100,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m010010_0	),
Adb51011100101	(	adb51011100101,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m010010_0	),
Adb51011100110	(	adb51011100110,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m010010_0	),
Adb51011100111	(	adb51011100111,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m010010_0	),
Adb51011101000	(	adb51011101000,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m010010_0	),
Adb51011101001	(	adb51011101001,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m010010_0	),
Adb51011101010	(	adb51011101010,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m010010_0	),
Adb51011101011	(	adb51011101011,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m010010_0	),
Adb51011101100	(	adb51011101100,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m010010_0	),
Adb51011101101	(	adb51011101101,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m010010_0	),
Adb51011101110	(	adb51011101110,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m010010_0	),
Adb51011101111	(	adb51011101111,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m010010_0	),
Adb51011110000	(	adb51011110000,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m010010_0	),
Adb51011110001	(	adb51011110001,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m010010_0	),
Adb51011110010	(	adb51011110010,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m010010_0	),
Adb51011110011	(	adb51011110011,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m010010_0	),
Adb51011110100	(	adb51011110100,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m010010_0	),
Adb51011110101	(	adb51011110101,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m010010_0	),
Adb51011110110	(	adb51011110110,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m010010_0	),
Adb51011110111	(	adb51011110111,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m010010_0	),
Adb51011111000	(	adb51011111000,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m010010_0	),
Adb51011111001	(	adb51011111001,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m010010_0	),
Adb51011111010	(	adb51011111010,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m010010_0	),
Adb51011111011	(	adb51011111011,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m010010_0	),
Adb51011111100	(	adb51011111100,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m010010_0	),
Adb51011111101	(	adb51011111101,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m010010_0	),
Adb51011111110	(	adb51011111110,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m010010_0	),
Adb51011111111	(	adb51011111111,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m010010_0	),
Adb51100000000	(	adb51100000000,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m001010_0	),
Adb51100000001	(	adb51100000001,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m001010_0	),
Adb51100000010	(	adb51100000010,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m001010_0	),
Adb51100000011	(	adb51100000011,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m001010_0	),
Adb51100000100	(	adb51100000100,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m001010_0	),
Adb51100000101	(	adb51100000101,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m001010_0	),
Adb51100000110	(	adb51100000110,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m001010_0	),
Adb51100000111	(	adb51100000111,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m001010_0	),
Adb51100001000	(	adb51100001000,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m001010_0	),
Adb51100001001	(	adb51100001001,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m001010_0	),
Adb51100001010	(	adb51100001010,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m001010_0	),
Adb51100001011	(	adb51100001011,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m001010_0	),
Adb51100001100	(	adb51100001100,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m001010_0	),
Adb51100001101	(	adb51100001101,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m001010_0	),
Adb51100001110	(	adb51100001110,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m001010_0	),
Adb51100001111	(	adb51100001111,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m001010_0	),
Adb51100010000	(	adb51100010000,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m001010_0	),
Adb51100010001	(	adb51100010001,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m001010_0	),
Adb51100010010	(	adb51100010010,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m001010_0	),
Adb51100010011	(	adb51100010011,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m001010_0	),
Adb51100010100	(	adb51100010100,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m001010_0	),
Adb51100010101	(	adb51100010101,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m001010_0	),
Adb51100010110	(	adb51100010110,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m001010_0	),
Adb51100010111	(	adb51100010111,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m001010_0	),
Adb51100011000	(	adb51100011000,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m001010_0	),
Adb51100011001	(	adb51100011001,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m001010_0	),
Adb51100011010	(	adb51100011010,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m001010_0	),
Adb51100011011	(	adb51100011011,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m001010_0	),
Adb51100011100	(	adb51100011100,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m001010_0	),
Adb51100011101	(	adb51100011101,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m001010_0	),
Adb51100011110	(	adb51100011110,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m001010_0	),
Adb51100011111	(	adb51100011111,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m001010_0	),
Adb51100100000	(	adb51100100000,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m001010_0	),
Adb51100100001	(	adb51100100001,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m001010_0	),
Adb51100100010	(	adb51100100010,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m001010_0	),
Adb51100100011	(	adb51100100011,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m001010_0	),
Adb51100100100	(	adb51100100100,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m001010_0	),
Adb51100100101	(	adb51100100101,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m001010_0	),
Adb51100100110	(	adb51100100110,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m001010_0	),
Adb51100100111	(	adb51100100111,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m001010_0	),
Adb51100101000	(	adb51100101000,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m001010_0	),
Adb51100101001	(	adb51100101001,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m001010_0	),
Adb51100101010	(	adb51100101010,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m001010_0	),
Adb51100101011	(	adb51100101011,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m001010_0	),
Adb51100101100	(	adb51100101100,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m001010_0	),
Adb51100101101	(	adb51100101101,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m001010_0	),
Adb51100101110	(	adb51100101110,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m001010_0	),
Adb51100101111	(	adb51100101111,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m001010_0	),
Adb51100110000	(	adb51100110000,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m001010_0	),
Adb51100110001	(	adb51100110001,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m001010_0	),
Adb51100110010	(	adb51100110010,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m001010_0	),
Adb51100110011	(	adb51100110011,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m001010_0	),
Adb51100110100	(	adb51100110100,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m001010_0	),
Adb51100110101	(	adb51100110101,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m001010_0	),
Adb51100110110	(	adb51100110110,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m001010_0	),
Adb51100110111	(	adb51100110111,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m001010_0	),
Adb51100111000	(	adb51100111000,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m001010_0	),
Adb51100111001	(	adb51100111001,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m001010_0	),
Adb51100111010	(	adb51100111010,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m001010_0	),
Adb51100111011	(	adb51100111011,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m001010_0	),
Adb51100111100	(	adb51100111100,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m001010_0	),
Adb51100111101	(	adb51100111101,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m001010_0	),
Adb51100111110	(	adb51100111110,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m001010_0	),
Adb51100111111	(	adb51100111111,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m001010_0	),
Adb51101000000	(	adb51101000000,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m001010_0	),
Adb51101000001	(	adb51101000001,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m001010_0	),
Adb51101000010	(	adb51101000010,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m001010_0	),
Adb51101000011	(	adb51101000011,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m001010_0	),
Adb51101000100	(	adb51101000100,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m001010_0	),
Adb51101000101	(	adb51101000101,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m001010_0	),
Adb51101000110	(	adb51101000110,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m001010_0	),
Adb51101000111	(	adb51101000111,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m001010_0	),
Adb51101001000	(	adb51101001000,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m001010_0	),
Adb51101001001	(	adb51101001001,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m001010_0	),
Adb51101001010	(	adb51101001010,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m001010_0	),
Adb51101001011	(	adb51101001011,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m001010_0	),
Adb51101001100	(	adb51101001100,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m001010_0	),
Adb51101001101	(	adb51101001101,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m001010_0	),
Adb51101001110	(	adb51101001110,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m001010_0	),
Adb51101001111	(	adb51101001111,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m001010_0	),
Adb51101010000	(	adb51101010000,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m001010_0	),
Adb51101010001	(	adb51101010001,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m001010_0	),
Adb51101010010	(	adb51101010010,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m001010_0	),
Adb51101010011	(	adb51101010011,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m001010_0	),
Adb51101010100	(	adb51101010100,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m001010_0	),
Adb51101010101	(	adb51101010101,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m001010_0	),
Adb51101010110	(	adb51101010110,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m001010_0	),
Adb51101010111	(	adb51101010111,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m001010_0	),
Adb51101011000	(	adb51101011000,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m001010_0	),
Adb51101011001	(	adb51101011001,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m001010_0	),
Adb51101011010	(	adb51101011010,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m001010_0	),
Adb51101011011	(	adb51101011011,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m001010_0	),
Adb51101011100	(	adb51101011100,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m001010_0	),
Adb51101011101	(	adb51101011101,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m001010_0	),
Adb51101011110	(	adb51101011110,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m001010_0	),
Adb51101011111	(	adb51101011111,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m001010_0	),
Adb51101100000	(	adb51101100000,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m001010_0	),
Adb51101100001	(	adb51101100001,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m001010_0	),
Adb51101100010	(	adb51101100010,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m001010_0	),
Adb51101100011	(	adb51101100011,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m001010_0	),
Adb51101100100	(	adb51101100100,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m001010_0	),
Adb51101100101	(	adb51101100101,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m001010_0	),
Adb51101100110	(	adb51101100110,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m001010_0	),
Adb51101100111	(	adb51101100111,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m001010_0	),
Adb51101101000	(	adb51101101000,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m001010_0	),
Adb51101101001	(	adb51101101001,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m001010_0	),
Adb51101101010	(	adb51101101010,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m001010_0	),
Adb51101101011	(	adb51101101011,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m001010_0	),
Adb51101101100	(	adb51101101100,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m001010_0	),
Adb51101101101	(	adb51101101101,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m001010_0	),
Adb51101101110	(	adb51101101110,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m001010_0	),
Adb51101101111	(	adb51101101111,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m001010_0	),
Adb51101110000	(	adb51101110000,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m001010_0	),
Adb51101110001	(	adb51101110001,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m001010_0	),
Adb51101110010	(	adb51101110010,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m001010_0	),
Adb51101110011	(	adb51101110011,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m001010_0	),
Adb51101110100	(	adb51101110100,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m001010_0	),
Adb51101110101	(	adb51101110101,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m001010_0	),
Adb51101110110	(	adb51101110110,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m001010_0	),
Adb51101110111	(	adb51101110111,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m001010_0	),
Adb51101111000	(	adb51101111000,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m001010_0	),
Adb51101111001	(	adb51101111001,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m001010_0	),
Adb51101111010	(	adb51101111010,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m001010_0	),
Adb51101111011	(	adb51101111011,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m001010_0	),
Adb51101111100	(	adb51101111100,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m001010_0	),
Adb51101111101	(	adb51101111101,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m001010_0	),
Adb51101111110	(	adb51101111110,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m001010_0	),
Adb51101111111	(	adb51101111111,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m001010_0	),
Adb51110000000	(	adb51110000000,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m000010_0	),
Adb51110000001	(	adb51110000001,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m000010_0	),
Adb51110000010	(	adb51110000010,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m000010_0	),
Adb51110000011	(	adb51110000011,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m000010_0	),
Adb51110000100	(	adb51110000100,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m000010_0	),
Adb51110000101	(	adb51110000101,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m000010_0	),
Adb51110000110	(	adb51110000110,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m000010_0	),
Adb51110000111	(	adb51110000111,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m000010_0	),
Adb51110001000	(	adb51110001000,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m000010_0	),
Adb51110001001	(	adb51110001001,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m000010_0	),
Adb51110001010	(	adb51110001010,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m000010_0	),
Adb51110001011	(	adb51110001011,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m000010_0	),
Adb51110001100	(	adb51110001100,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m000010_0	),
Adb51110001101	(	adb51110001101,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m000010_0	),
Adb51110001110	(	adb51110001110,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m000010_0	),
Adb51110001111	(	adb51110001111,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m000010_0	),
Adb51110010000	(	adb51110010000,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m000010_0	),
Adb51110010001	(	adb51110010001,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m000010_0	),
Adb51110010010	(	adb51110010010,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m000010_0	),
Adb51110010011	(	adb51110010011,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m000010_0	),
Adb51110010100	(	adb51110010100,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m000010_0	),
Adb51110010101	(	adb51110010101,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m000010_0	),
Adb51110010110	(	adb51110010110,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m000010_0	),
Adb51110010111	(	adb51110010111,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m000010_0	),
Adb51110011000	(	adb51110011000,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m000010_0	),
Adb51110011001	(	adb51110011001,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m000010_0	),
Adb51110011010	(	adb51110011010,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m000010_0	),
Adb51110011011	(	adb51110011011,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m000010_0	),
Adb51110011100	(	adb51110011100,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m000010_0	),
Adb51110011101	(	adb51110011101,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m000010_0	),
Adb51110011110	(	adb51110011110,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m000010_0	),
Adb51110011111	(	adb51110011111,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m000010_0	),
Adb51110100000	(	adb51110100000,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m000010_0	),
Adb51110100001	(	adb51110100001,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m000010_0	),
Adb51110100010	(	adb51110100010,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m000010_0	),
Adb51110100011	(	adb51110100011,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m000010_0	),
Adb51110100100	(	adb51110100100,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m000010_0	),
Adb51110100101	(	adb51110100101,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m000010_0	),
Adb51110100110	(	adb51110100110,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m000010_0	),
Adb51110100111	(	adb51110100111,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m000010_0	),
Adb51110101000	(	adb51110101000,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m000010_0	),
Adb51110101001	(	adb51110101001,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m000010_0	),
Adb51110101010	(	adb51110101010,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m000010_0	),
Adb51110101011	(	adb51110101011,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m000010_0	),
Adb51110101100	(	adb51110101100,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m000010_0	),
Adb51110101101	(	adb51110101101,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m000010_0	),
Adb51110101110	(	adb51110101110,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m000010_0	),
Adb51110101111	(	adb51110101111,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m000010_0	),
Adb51110110000	(	adb51110110000,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m000010_0	),
Adb51110110001	(	adb51110110001,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m000010_0	),
Adb51110110010	(	adb51110110010,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m000010_0	),
Adb51110110011	(	adb51110110011,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m000010_0	),
Adb51110110100	(	adb51110110100,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m000010_0	),
Adb51110110101	(	adb51110110101,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m000010_0	),
Adb51110110110	(	adb51110110110,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m000010_0	),
Adb51110110111	(	adb51110110111,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m000010_0	),
Adb51110111000	(	adb51110111000,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m000010_0	),
Adb51110111001	(	adb51110111001,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m000010_0	),
Adb51110111010	(	adb51110111010,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m000010_0	),
Adb51110111011	(	adb51110111011,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m000010_0	),
Adb51110111100	(	adb51110111100,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m000010_0	),
Adb51110111101	(	adb51110111101,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m000010_0	),
Adb51110111110	(	adb51110111110,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m000010_0	),
Adb51110111111	(	adb51110111111,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m000010_0	),
Adb51111000000	(	adb51111000000,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m000010_0	),
Adb51111000001	(	adb51111000001,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m000010_0	),
Adb51111000010	(	adb51111000010,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m000010_0	),
Adb51111000011	(	adb51111000011,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m000010_0	),
Adb51111000100	(	adb51111000100,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m000010_0	),
Adb51111000101	(	adb51111000101,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m000010_0	),
Adb51111000110	(	adb51111000110,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m000010_0	),
Adb51111000111	(	adb51111000111,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m000010_0	),
Adb51111001000	(	adb51111001000,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m000010_0	),
Adb51111001001	(	adb51111001001,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m000010_0	),
Adb51111001010	(	adb51111001010,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m000010_0	),
Adb51111001011	(	adb51111001011,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m000010_0	),
Adb51111001100	(	adb51111001100,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m000010_0	),
Adb51111001101	(	adb51111001101,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m000010_0	),
Adb51111001110	(	adb51111001110,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m000010_0	),
Adb51111001111	(	adb51111001111,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m000010_0	),
Adb51111010000	(	adb51111010000,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m000010_0	),
Adb51111010001	(	adb51111010001,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m000010_0	),
Adb51111010010	(	adb51111010010,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m000010_0	),
Adb51111010011	(	adb51111010011,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m000010_0	),
Adb51111010100	(	adb51111010100,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m000010_0	),
Adb51111010101	(	adb51111010101,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m000010_0	),
Adb51111010110	(	adb51111010110,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m000010_0	),
Adb51111010111	(	adb51111010111,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m000010_0	),
Adb51111011000	(	adb51111011000,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m000010_0	),
Adb51111011001	(	adb51111011001,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m000010_0	),
Adb51111011010	(	adb51111011010,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m000010_0	),
Adb51111011011	(	adb51111011011,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m000010_0	),
Adb51111011100	(	adb51111011100,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m000010_0	),
Adb51111011101	(	adb51111011101,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m000010_0	),
Adb51111011110	(	adb51111011110,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m000010_0	),
Adb51111011111	(	adb51111011111,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m000010_0	),
Adb51111100000	(	adb51111100000,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m000010_0	),
Adb51111100001	(	adb51111100001,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m000010_0	),
Adb51111100010	(	adb51111100010,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m000010_0	),
Adb51111100011	(	adb51111100011,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m000010_0	),
Adb51111100100	(	adb51111100100,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m000010_0	),
Adb51111100101	(	adb51111100101,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m000010_0	),
Adb51111100110	(	adb51111100110,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m000010_0	),
Adb51111100111	(	adb51111100111,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m000010_0	),
Adb51111101000	(	adb51111101000,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m000010_0	),
Adb51111101001	(	adb51111101001,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m000010_0	),
Adb51111101010	(	adb51111101010,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m000010_0	),
Adb51111101011	(	adb51111101011,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m000010_0	),
Adb51111101100	(	adb51111101100,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m000010_0	),
Adb51111101101	(	adb51111101101,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m000010_0	),
Adb51111101110	(	adb51111101110,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m000010_0	),
Adb51111101111	(	adb51111101111,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m000010_0	),
Adb51111110000	(	adb51111110000,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m000010_0	),
Adb51111110001	(	adb51111110001,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m000010_0	),
Adb51111110010	(	adb51111110010,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m000010_0	),
Adb51111110011	(	adb51111110011,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m000010_0	),
Adb51111110100	(	adb51111110100,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m000010_0	),
Adb51111110101	(	adb51111110101,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m000010_0	),
Adb51111110110	(	adb51111110110,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m000010_0	),
Adb51111110111	(	adb51111110111,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m000010_0	),
Adb51111111000	(	adb51111111000,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m000010_0	),
Adb51111111001	(	adb51111111001,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m000010_0	),
Adb51111111010	(	adb51111111010,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m000010_0	),
Adb51111111011	(	adb51111111011,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m000010_0	),
Adb51111111100	(	adb51111111100,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m000010_0	),
Adb51111111101	(	adb51111111101,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m000010_0	),
Adb51111111110	(	adb51111111110,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m000010_0	),
Adb51111111111	(	adb51111111111,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m000010_0	),
       Adb600(adb600,n0011,n0010,n0009,m0009),
       Adb601(adb601,n0011,n0010,m0009,m0009),
       Adb610(adb610,n0011,m0010,n0009,m0009),
       Adb611(adb611,n0011,m0010,m0009,m0009),
Adb60000000000	(	adb60000000000,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m111001_0	),
Adb60000000001	(	adb60000000001,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m111001_0	),
Adb60000000010	(	adb60000000010,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m111001_0	),
Adb60000000011	(	adb60000000011,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m111001_0	),
Adb60000000100	(	adb60000000100,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m111001_0	),
Adb60000000101	(	adb60000000101,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m111001_0	),
Adb60000000110	(	adb60000000110,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m111001_0	),
Adb60000000111	(	adb60000000111,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m111001_0	),
Adb60000001000	(	adb60000001000,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m111001_0	),
Adb60000001001	(	adb60000001001,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m111001_0	),
Adb60000001010	(	adb60000001010,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m111001_0	),
Adb60000001011	(	adb60000001011,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m111001_0	),
Adb60000001100	(	adb60000001100,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m111001_0	),
Adb60000001101	(	adb60000001101,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m111001_0	),
Adb60000001110	(	adb60000001110,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m111001_0	),
Adb60000001111	(	adb60000001111,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m111001_0	),
Adb60000010000	(	adb60000010000,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m111001_0	),
Adb60000010001	(	adb60000010001,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m111001_0	),
Adb60000010010	(	adb60000010010,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m111001_0	),
Adb60000010011	(	adb60000010011,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m111001_0	),
Adb60000010100	(	adb60000010100,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m111001_0	),
Adb60000010101	(	adb60000010101,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m111001_0	),
Adb60000010110	(	adb60000010110,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m111001_0	),
Adb60000010111	(	adb60000010111,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m111001_0	),
Adb60000011000	(	adb60000011000,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m111001_0	),
Adb60000011001	(	adb60000011001,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m111001_0	),
Adb60000011010	(	adb60000011010,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m111001_0	),
Adb60000011011	(	adb60000011011,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m111001_0	),
Adb60000011100	(	adb60000011100,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m111001_0	),
Adb60000011101	(	adb60000011101,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m111001_0	),
Adb60000011110	(	adb60000011110,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m111001_0	),
Adb60000011111	(	adb60000011111,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m111001_0	),
Adb60000100000	(	adb60000100000,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m111001_0	),
Adb60000100001	(	adb60000100001,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m111001_0	),
Adb60000100010	(	adb60000100010,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m111001_0	),
Adb60000100011	(	adb60000100011,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m111001_0	),
Adb60000100100	(	adb60000100100,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m111001_0	),
Adb60000100101	(	adb60000100101,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m111001_0	),
Adb60000100110	(	adb60000100110,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m111001_0	),
Adb60000100111	(	adb60000100111,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m111001_0	),
Adb60000101000	(	adb60000101000,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m111001_0	),
Adb60000101001	(	adb60000101001,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m111001_0	),
Adb60000101010	(	adb60000101010,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m111001_0	),
Adb60000101011	(	adb60000101011,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m111001_0	),
Adb60000101100	(	adb60000101100,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m111001_0	),
Adb60000101101	(	adb60000101101,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m111001_0	),
Adb60000101110	(	adb60000101110,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m111001_0	),
Adb60000101111	(	adb60000101111,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m111001_0	),
Adb60000110000	(	adb60000110000,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m111001_0	),
Adb60000110001	(	adb60000110001,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m111001_0	),
Adb60000110010	(	adb60000110010,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m111001_0	),
Adb60000110011	(	adb60000110011,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m111001_0	),
Adb60000110100	(	adb60000110100,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m111001_0	),
Adb60000110101	(	adb60000110101,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m111001_0	),
Adb60000110110	(	adb60000110110,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m111001_0	),
Adb60000110111	(	adb60000110111,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m111001_0	),
Adb60000111000	(	adb60000111000,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m111001_0	),
Adb60000111001	(	adb60000111001,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m111001_0	),
Adb60000111010	(	adb60000111010,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m111001_0	),
Adb60000111011	(	adb60000111011,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m111001_0	),
Adb60000111100	(	adb60000111100,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m111001_0	),
Adb60000111101	(	adb60000111101,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m111001_0	),
Adb60000111110	(	adb60000111110,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m111001_0	),
Adb60000111111	(	adb60000111111,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m111001_0	),
Adb60001000000	(	adb60001000000,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m111001_0	),
Adb60001000001	(	adb60001000001,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m111001_0	),
Adb60001000010	(	adb60001000010,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m111001_0	),
Adb60001000011	(	adb60001000011,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m111001_0	),
Adb60001000100	(	adb60001000100,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m111001_0	),
Adb60001000101	(	adb60001000101,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m111001_0	),
Adb60001000110	(	adb60001000110,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m111001_0	),
Adb60001000111	(	adb60001000111,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m111001_0	),
Adb60001001000	(	adb60001001000,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m111001_0	),
Adb60001001001	(	adb60001001001,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m111001_0	),
Adb60001001010	(	adb60001001010,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m111001_0	),
Adb60001001011	(	adb60001001011,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m111001_0	),
Adb60001001100	(	adb60001001100,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m111001_0	),
Adb60001001101	(	adb60001001101,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m111001_0	),
Adb60001001110	(	adb60001001110,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m111001_0	),
Adb60001001111	(	adb60001001111,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m111001_0	),
Adb60001010000	(	adb60001010000,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m111001_0	),
Adb60001010001	(	adb60001010001,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m111001_0	),
Adb60001010010	(	adb60001010010,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m111001_0	),
Adb60001010011	(	adb60001010011,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m111001_0	),
Adb60001010100	(	adb60001010100,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m111001_0	),
Adb60001010101	(	adb60001010101,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m111001_0	),
Adb60001010110	(	adb60001010110,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m111001_0	),
Adb60001010111	(	adb60001010111,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m111001_0	),
Adb60001011000	(	adb60001011000,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m111001_0	),
Adb60001011001	(	adb60001011001,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m111001_0	),
Adb60001011010	(	adb60001011010,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m111001_0	),
Adb60001011011	(	adb60001011011,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m111001_0	),
Adb60001011100	(	adb60001011100,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m111001_0	),
Adb60001011101	(	adb60001011101,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m111001_0	),
Adb60001011110	(	adb60001011110,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m111001_0	),
Adb60001011111	(	adb60001011111,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m111001_0	),
Adb60001100000	(	adb60001100000,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m111001_0	),
Adb60001100001	(	adb60001100001,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m111001_0	),
Adb60001100010	(	adb60001100010,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m111001_0	),
Adb60001100011	(	adb60001100011,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m111001_0	),
Adb60001100100	(	adb60001100100,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m111001_0	),
Adb60001100101	(	adb60001100101,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m111001_0	),
Adb60001100110	(	adb60001100110,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m111001_0	),
Adb60001100111	(	adb60001100111,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m111001_0	),
Adb60001101000	(	adb60001101000,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m111001_0	),
Adb60001101001	(	adb60001101001,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m111001_0	),
Adb60001101010	(	adb60001101010,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m111001_0	),
Adb60001101011	(	adb60001101011,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m111001_0	),
Adb60001101100	(	adb60001101100,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m111001_0	),
Adb60001101101	(	adb60001101101,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m111001_0	),
Adb60001101110	(	adb60001101110,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m111001_0	),
Adb60001101111	(	adb60001101111,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m111001_0	),
Adb60001110000	(	adb60001110000,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m111001_0	),
Adb60001110001	(	adb60001110001,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m111001_0	),
Adb60001110010	(	adb60001110010,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m111001_0	),
Adb60001110011	(	adb60001110011,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m111001_0	),
Adb60001110100	(	adb60001110100,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m111001_0	),
Adb60001110101	(	adb60001110101,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m111001_0	),
Adb60001110110	(	adb60001110110,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m111001_0	),
Adb60001110111	(	adb60001110111,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m111001_0	),
Adb60001111000	(	adb60001111000,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m111001_0	),
Adb60001111001	(	adb60001111001,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m111001_0	),
Adb60001111010	(	adb60001111010,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m111001_0	),
Adb60001111011	(	adb60001111011,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m111001_0	),
Adb60001111100	(	adb60001111100,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m111001_0	),
Adb60001111101	(	adb60001111101,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m111001_0	),
Adb60001111110	(	adb60001111110,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m111001_0	),
Adb60001111111	(	adb60001111111,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m111001_0	),
Adb60010000000	(	adb60010000000,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m110001_0	),
Adb60010000001	(	adb60010000001,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m110001_0	),
Adb60010000010	(	adb60010000010,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m110001_0	),
Adb60010000011	(	adb60010000011,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m110001_0	),
Adb60010000100	(	adb60010000100,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m110001_0	),
Adb60010000101	(	adb60010000101,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m110001_0	),
Adb60010000110	(	adb60010000110,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m110001_0	),
Adb60010000111	(	adb60010000111,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m110001_0	),
Adb60010001000	(	adb60010001000,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m110001_0	),
Adb60010001001	(	adb60010001001,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m110001_0	),
Adb60010001010	(	adb60010001010,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m110001_0	),
Adb60010001011	(	adb60010001011,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m110001_0	),
Adb60010001100	(	adb60010001100,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m110001_0	),
Adb60010001101	(	adb60010001101,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m110001_0	),
Adb60010001110	(	adb60010001110,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m110001_0	),
Adb60010001111	(	adb60010001111,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m110001_0	),
Adb60010010000	(	adb60010010000,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m110001_0	),
Adb60010010001	(	adb60010010001,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m110001_0	),
Adb60010010010	(	adb60010010010,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m110001_0	),
Adb60010010011	(	adb60010010011,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m110001_0	),
Adb60010010100	(	adb60010010100,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m110001_0	),
Adb60010010101	(	adb60010010101,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m110001_0	),
Adb60010010110	(	adb60010010110,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m110001_0	),
Adb60010010111	(	adb60010010111,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m110001_0	),
Adb60010011000	(	adb60010011000,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m110001_0	),
Adb60010011001	(	adb60010011001,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m110001_0	),
Adb60010011010	(	adb60010011010,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m110001_0	),
Adb60010011011	(	adb60010011011,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m110001_0	),
Adb60010011100	(	adb60010011100,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m110001_0	),
Adb60010011101	(	adb60010011101,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m110001_0	),
Adb60010011110	(	adb60010011110,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m110001_0	),
Adb60010011111	(	adb60010011111,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m110001_0	),
Adb60010100000	(	adb60010100000,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m110001_0	),
Adb60010100001	(	adb60010100001,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m110001_0	),
Adb60010100010	(	adb60010100010,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m110001_0	),
Adb60010100011	(	adb60010100011,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m110001_0	),
Adb60010100100	(	adb60010100100,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m110001_0	),
Adb60010100101	(	adb60010100101,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m110001_0	),
Adb60010100110	(	adb60010100110,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m110001_0	),
Adb60010100111	(	adb60010100111,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m110001_0	),
Adb60010101000	(	adb60010101000,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m110001_0	),
Adb60010101001	(	adb60010101001,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m110001_0	),
Adb60010101010	(	adb60010101010,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m110001_0	),
Adb60010101011	(	adb60010101011,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m110001_0	),
Adb60010101100	(	adb60010101100,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m110001_0	),
Adb60010101101	(	adb60010101101,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m110001_0	),
Adb60010101110	(	adb60010101110,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m110001_0	),
Adb60010101111	(	adb60010101111,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m110001_0	),
Adb60010110000	(	adb60010110000,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m110001_0	),
Adb60010110001	(	adb60010110001,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m110001_0	),
Adb60010110010	(	adb60010110010,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m110001_0	),
Adb60010110011	(	adb60010110011,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m110001_0	),
Adb60010110100	(	adb60010110100,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m110001_0	),
Adb60010110101	(	adb60010110101,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m110001_0	),
Adb60010110110	(	adb60010110110,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m110001_0	),
Adb60010110111	(	adb60010110111,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m110001_0	),
Adb60010111000	(	adb60010111000,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m110001_0	),
Adb60010111001	(	adb60010111001,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m110001_0	),
Adb60010111010	(	adb60010111010,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m110001_0	),
Adb60010111011	(	adb60010111011,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m110001_0	),
Adb60010111100	(	adb60010111100,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m110001_0	),
Adb60010111101	(	adb60010111101,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m110001_0	),
Adb60010111110	(	adb60010111110,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m110001_0	),
Adb60010111111	(	adb60010111111,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m110001_0	),
Adb60011000000	(	adb60011000000,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m110001_0	),
Adb60011000001	(	adb60011000001,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m110001_0	),
Adb60011000010	(	adb60011000010,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m110001_0	),
Adb60011000011	(	adb60011000011,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m110001_0	),
Adb60011000100	(	adb60011000100,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m110001_0	),
Adb60011000101	(	adb60011000101,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m110001_0	),
Adb60011000110	(	adb60011000110,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m110001_0	),
Adb60011000111	(	adb60011000111,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m110001_0	),
Adb60011001000	(	adb60011001000,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m110001_0	),
Adb60011001001	(	adb60011001001,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m110001_0	),
Adb60011001010	(	adb60011001010,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m110001_0	),
Adb60011001011	(	adb60011001011,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m110001_0	),
Adb60011001100	(	adb60011001100,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m110001_0	),
Adb60011001101	(	adb60011001101,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m110001_0	),
Adb60011001110	(	adb60011001110,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m110001_0	),
Adb60011001111	(	adb60011001111,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m110001_0	),
Adb60011010000	(	adb60011010000,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m110001_0	),
Adb60011010001	(	adb60011010001,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m110001_0	),
Adb60011010010	(	adb60011010010,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m110001_0	),
Adb60011010011	(	adb60011010011,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m110001_0	),
Adb60011010100	(	adb60011010100,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m110001_0	),
Adb60011010101	(	adb60011010101,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m110001_0	),
Adb60011010110	(	adb60011010110,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m110001_0	),
Adb60011010111	(	adb60011010111,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m110001_0	),
Adb60011011000	(	adb60011011000,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m110001_0	),
Adb60011011001	(	adb60011011001,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m110001_0	),
Adb60011011010	(	adb60011011010,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m110001_0	),
Adb60011011011	(	adb60011011011,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m110001_0	),
Adb60011011100	(	adb60011011100,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m110001_0	),
Adb60011011101	(	adb60011011101,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m110001_0	),
Adb60011011110	(	adb60011011110,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m110001_0	),
Adb60011011111	(	adb60011011111,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m110001_0	),
Adb60011100000	(	adb60011100000,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m110001_0	),
Adb60011100001	(	adb60011100001,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m110001_0	),
Adb60011100010	(	adb60011100010,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m110001_0	),
Adb60011100011	(	adb60011100011,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m110001_0	),
Adb60011100100	(	adb60011100100,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m110001_0	),
Adb60011100101	(	adb60011100101,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m110001_0	),
Adb60011100110	(	adb60011100110,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m110001_0	),
Adb60011100111	(	adb60011100111,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m110001_0	),
Adb60011101000	(	adb60011101000,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m110001_0	),
Adb60011101001	(	adb60011101001,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m110001_0	),
Adb60011101010	(	adb60011101010,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m110001_0	),
Adb60011101011	(	adb60011101011,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m110001_0	),
Adb60011101100	(	adb60011101100,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m110001_0	),
Adb60011101101	(	adb60011101101,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m110001_0	),
Adb60011101110	(	adb60011101110,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m110001_0	),
Adb60011101111	(	adb60011101111,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m110001_0	),
Adb60011110000	(	adb60011110000,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m110001_0	),
Adb60011110001	(	adb60011110001,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m110001_0	),
Adb60011110010	(	adb60011110010,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m110001_0	),
Adb60011110011	(	adb60011110011,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m110001_0	),
Adb60011110100	(	adb60011110100,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m110001_0	),
Adb60011110101	(	adb60011110101,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m110001_0	),
Adb60011110110	(	adb60011110110,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m110001_0	),
Adb60011110111	(	adb60011110111,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m110001_0	),
Adb60011111000	(	adb60011111000,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m110001_0	),
Adb60011111001	(	adb60011111001,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m110001_0	),
Adb60011111010	(	adb60011111010,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m110001_0	),
Adb60011111011	(	adb60011111011,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m110001_0	),
Adb60011111100	(	adb60011111100,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m110001_0	),
Adb60011111101	(	adb60011111101,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m110001_0	),
Adb60011111110	(	adb60011111110,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m110001_0	),
Adb60011111111	(	adb60011111111,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m110001_0	),
Adb60100000000	(	adb60100000000,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m101001_0	),
Adb60100000001	(	adb60100000001,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m101001_0	),
Adb60100000010	(	adb60100000010,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m101001_0	),
Adb60100000011	(	adb60100000011,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m101001_0	),
Adb60100000100	(	adb60100000100,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m101001_0	),
Adb60100000101	(	adb60100000101,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m101001_0	),
Adb60100000110	(	adb60100000110,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m101001_0	),
Adb60100000111	(	adb60100000111,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m101001_0	),
Adb60100001000	(	adb60100001000,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m101001_0	),
Adb60100001001	(	adb60100001001,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m101001_0	),
Adb60100001010	(	adb60100001010,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m101001_0	),
Adb60100001011	(	adb60100001011,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m101001_0	),
Adb60100001100	(	adb60100001100,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m101001_0	),
Adb60100001101	(	adb60100001101,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m101001_0	),
Adb60100001110	(	adb60100001110,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m101001_0	),
Adb60100001111	(	adb60100001111,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m101001_0	),
Adb60100010000	(	adb60100010000,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m101001_0	),
Adb60100010001	(	adb60100010001,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m101001_0	),
Adb60100010010	(	adb60100010010,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m101001_0	),
Adb60100010011	(	adb60100010011,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m101001_0	),
Adb60100010100	(	adb60100010100,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m101001_0	),
Adb60100010101	(	adb60100010101,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m101001_0	),
Adb60100010110	(	adb60100010110,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m101001_0	),
Adb60100010111	(	adb60100010111,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m101001_0	),
Adb60100011000	(	adb60100011000,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m101001_0	),
Adb60100011001	(	adb60100011001,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m101001_0	),
Adb60100011010	(	adb60100011010,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m101001_0	),
Adb60100011011	(	adb60100011011,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m101001_0	),
Adb60100011100	(	adb60100011100,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m101001_0	),
Adb60100011101	(	adb60100011101,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m101001_0	),
Adb60100011110	(	adb60100011110,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m101001_0	),
Adb60100011111	(	adb60100011111,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m101001_0	),
Adb60100100000	(	adb60100100000,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m101001_0	),
Adb60100100001	(	adb60100100001,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m101001_0	),
Adb60100100010	(	adb60100100010,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m101001_0	),
Adb60100100011	(	adb60100100011,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m101001_0	),
Adb60100100100	(	adb60100100100,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m101001_0	),
Adb60100100101	(	adb60100100101,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m101001_0	),
Adb60100100110	(	adb60100100110,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m101001_0	),
Adb60100100111	(	adb60100100111,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m101001_0	),
Adb60100101000	(	adb60100101000,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m101001_0	),
Adb60100101001	(	adb60100101001,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m101001_0	),
Adb60100101010	(	adb60100101010,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m101001_0	),
Adb60100101011	(	adb60100101011,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m101001_0	),
Adb60100101100	(	adb60100101100,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m101001_0	),
Adb60100101101	(	adb60100101101,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m101001_0	),
Adb60100101110	(	adb60100101110,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m101001_0	),
Adb60100101111	(	adb60100101111,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m101001_0	),
Adb60100110000	(	adb60100110000,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m101001_0	),
Adb60100110001	(	adb60100110001,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m101001_0	),
Adb60100110010	(	adb60100110010,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m101001_0	),
Adb60100110011	(	adb60100110011,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m101001_0	),
Adb60100110100	(	adb60100110100,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m101001_0	),
Adb60100110101	(	adb60100110101,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m101001_0	),
Adb60100110110	(	adb60100110110,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m101001_0	),
Adb60100110111	(	adb60100110111,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m101001_0	),
Adb60100111000	(	adb60100111000,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m101001_0	),
Adb60100111001	(	adb60100111001,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m101001_0	),
Adb60100111010	(	adb60100111010,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m101001_0	),
Adb60100111011	(	adb60100111011,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m101001_0	),
Adb60100111100	(	adb60100111100,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m101001_0	),
Adb60100111101	(	adb60100111101,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m101001_0	),
Adb60100111110	(	adb60100111110,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m101001_0	),
Adb60100111111	(	adb60100111111,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m101001_0	),
Adb60101000000	(	adb60101000000,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m101001_0	),
Adb60101000001	(	adb60101000001,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m101001_0	),
Adb60101000010	(	adb60101000010,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m101001_0	),
Adb60101000011	(	adb60101000011,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m101001_0	),
Adb60101000100	(	adb60101000100,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m101001_0	),
Adb60101000101	(	adb60101000101,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m101001_0	),
Adb60101000110	(	adb60101000110,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m101001_0	),
Adb60101000111	(	adb60101000111,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m101001_0	),
Adb60101001000	(	adb60101001000,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m101001_0	),
Adb60101001001	(	adb60101001001,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m101001_0	),
Adb60101001010	(	adb60101001010,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m101001_0	),
Adb60101001011	(	adb60101001011,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m101001_0	),
Adb60101001100	(	adb60101001100,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m101001_0	),
Adb60101001101	(	adb60101001101,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m101001_0	),
Adb60101001110	(	adb60101001110,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m101001_0	),
Adb60101001111	(	adb60101001111,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m101001_0	),
Adb60101010000	(	adb60101010000,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m101001_0	),
Adb60101010001	(	adb60101010001,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m101001_0	),
Adb60101010010	(	adb60101010010,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m101001_0	),
Adb60101010011	(	adb60101010011,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m101001_0	),
Adb60101010100	(	adb60101010100,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m101001_0	),
Adb60101010101	(	adb60101010101,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m101001_0	),
Adb60101010110	(	adb60101010110,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m101001_0	),
Adb60101010111	(	adb60101010111,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m101001_0	),
Adb60101011000	(	adb60101011000,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m101001_0	),
Adb60101011001	(	adb60101011001,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m101001_0	),
Adb60101011010	(	adb60101011010,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m101001_0	),
Adb60101011011	(	adb60101011011,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m101001_0	),
Adb60101011100	(	adb60101011100,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m101001_0	),
Adb60101011101	(	adb60101011101,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m101001_0	),
Adb60101011110	(	adb60101011110,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m101001_0	),
Adb60101011111	(	adb60101011111,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m101001_0	),
Adb60101100000	(	adb60101100000,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m101001_0	),
Adb60101100001	(	adb60101100001,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m101001_0	),
Adb60101100010	(	adb60101100010,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m101001_0	),
Adb60101100011	(	adb60101100011,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m101001_0	),
Adb60101100100	(	adb60101100100,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m101001_0	),
Adb60101100101	(	adb60101100101,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m101001_0	),
Adb60101100110	(	adb60101100110,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m101001_0	),
Adb60101100111	(	adb60101100111,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m101001_0	),
Adb60101101000	(	adb60101101000,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m101001_0	),
Adb60101101001	(	adb60101101001,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m101001_0	),
Adb60101101010	(	adb60101101010,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m101001_0	),
Adb60101101011	(	adb60101101011,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m101001_0	),
Adb60101101100	(	adb60101101100,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m101001_0	),
Adb60101101101	(	adb60101101101,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m101001_0	),
Adb60101101110	(	adb60101101110,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m101001_0	),
Adb60101101111	(	adb60101101111,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m101001_0	),
Adb60101110000	(	adb60101110000,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m101001_0	),
Adb60101110001	(	adb60101110001,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m101001_0	),
Adb60101110010	(	adb60101110010,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m101001_0	),
Adb60101110011	(	adb60101110011,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m101001_0	),
Adb60101110100	(	adb60101110100,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m101001_0	),
Adb60101110101	(	adb60101110101,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m101001_0	),
Adb60101110110	(	adb60101110110,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m101001_0	),
Adb60101110111	(	adb60101110111,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m101001_0	),
Adb60101111000	(	adb60101111000,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m101001_0	),
Adb60101111001	(	adb60101111001,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m101001_0	),
Adb60101111010	(	adb60101111010,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m101001_0	),
Adb60101111011	(	adb60101111011,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m101001_0	),
Adb60101111100	(	adb60101111100,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m101001_0	),
Adb60101111101	(	adb60101111101,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m101001_0	),
Adb60101111110	(	adb60101111110,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m101001_0	),
Adb60101111111	(	adb60101111111,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m101001_0	),
Adb60110000000	(	adb60110000000,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m100001_0	),
Adb60110000001	(	adb60110000001,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m100001_0	),
Adb60110000010	(	adb60110000010,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m100001_0	),
Adb60110000011	(	adb60110000011,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m100001_0	),
Adb60110000100	(	adb60110000100,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m100001_0	),
Adb60110000101	(	adb60110000101,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m100001_0	),
Adb60110000110	(	adb60110000110,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m100001_0	),
Adb60110000111	(	adb60110000111,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m100001_0	),
Adb60110001000	(	adb60110001000,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m100001_0	),
Adb60110001001	(	adb60110001001,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m100001_0	),
Adb60110001010	(	adb60110001010,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m100001_0	),
Adb60110001011	(	adb60110001011,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m100001_0	),
Adb60110001100	(	adb60110001100,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m100001_0	),
Adb60110001101	(	adb60110001101,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m100001_0	),
Adb60110001110	(	adb60110001110,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m100001_0	),
Adb60110001111	(	adb60110001111,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m100001_0	),
Adb60110010000	(	adb60110010000,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m100001_0	),
Adb60110010001	(	adb60110010001,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m100001_0	),
Adb60110010010	(	adb60110010010,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m100001_0	),
Adb60110010011	(	adb60110010011,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m100001_0	),
Adb60110010100	(	adb60110010100,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m100001_0	),
Adb60110010101	(	adb60110010101,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m100001_0	),
Adb60110010110	(	adb60110010110,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m100001_0	),
Adb60110010111	(	adb60110010111,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m100001_0	),
Adb60110011000	(	adb60110011000,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m100001_0	),
Adb60110011001	(	adb60110011001,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m100001_0	),
Adb60110011010	(	adb60110011010,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m100001_0	),
Adb60110011011	(	adb60110011011,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m100001_0	),
Adb60110011100	(	adb60110011100,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m100001_0	),
Adb60110011101	(	adb60110011101,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m100001_0	),
Adb60110011110	(	adb60110011110,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m100001_0	),
Adb60110011111	(	adb60110011111,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m100001_0	),
Adb60110100000	(	adb60110100000,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m100001_0	),
Adb60110100001	(	adb60110100001,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m100001_0	),
Adb60110100010	(	adb60110100010,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m100001_0	),
Adb60110100011	(	adb60110100011,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m100001_0	),
Adb60110100100	(	adb60110100100,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m100001_0	),
Adb60110100101	(	adb60110100101,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m100001_0	),
Adb60110100110	(	adb60110100110,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m100001_0	),
Adb60110100111	(	adb60110100111,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m100001_0	),
Adb60110101000	(	adb60110101000,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m100001_0	),
Adb60110101001	(	adb60110101001,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m100001_0	),
Adb60110101010	(	adb60110101010,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m100001_0	),
Adb60110101011	(	adb60110101011,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m100001_0	),
Adb60110101100	(	adb60110101100,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m100001_0	),
Adb60110101101	(	adb60110101101,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m100001_0	),
Adb60110101110	(	adb60110101110,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m100001_0	),
Adb60110101111	(	adb60110101111,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m100001_0	),
Adb60110110000	(	adb60110110000,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m100001_0	),
Adb60110110001	(	adb60110110001,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m100001_0	),
Adb60110110010	(	adb60110110010,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m100001_0	),
Adb60110110011	(	adb60110110011,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m100001_0	),
Adb60110110100	(	adb60110110100,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m100001_0	),
Adb60110110101	(	adb60110110101,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m100001_0	),
Adb60110110110	(	adb60110110110,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m100001_0	),
Adb60110110111	(	adb60110110111,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m100001_0	),
Adb60110111000	(	adb60110111000,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m100001_0	),
Adb60110111001	(	adb60110111001,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m100001_0	),
Adb60110111010	(	adb60110111010,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m100001_0	),
Adb60110111011	(	adb60110111011,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m100001_0	),
Adb60110111100	(	adb60110111100,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m100001_0	),
Adb60110111101	(	adb60110111101,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m100001_0	),
Adb60110111110	(	adb60110111110,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m100001_0	),
Adb60110111111	(	adb60110111111,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m100001_0	),
Adb60111000000	(	adb60111000000,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m100001_0	),
Adb60111000001	(	adb60111000001,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m100001_0	),
Adb60111000010	(	adb60111000010,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m100001_0	),
Adb60111000011	(	adb60111000011,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m100001_0	),
Adb60111000100	(	adb60111000100,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m100001_0	),
Adb60111000101	(	adb60111000101,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m100001_0	),
Adb60111000110	(	adb60111000110,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m100001_0	),
Adb60111000111	(	adb60111000111,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m100001_0	),
Adb60111001000	(	adb60111001000,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m100001_0	),
Adb60111001001	(	adb60111001001,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m100001_0	),
Adb60111001010	(	adb60111001010,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m100001_0	),
Adb60111001011	(	adb60111001011,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m100001_0	),
Adb60111001100	(	adb60111001100,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m100001_0	),
Adb60111001101	(	adb60111001101,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m100001_0	),
Adb60111001110	(	adb60111001110,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m100001_0	),
Adb60111001111	(	adb60111001111,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m100001_0	),
Adb60111010000	(	adb60111010000,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m100001_0	),
Adb60111010001	(	adb60111010001,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m100001_0	),
Adb60111010010	(	adb60111010010,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m100001_0	),
Adb60111010011	(	adb60111010011,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m100001_0	),
Adb60111010100	(	adb60111010100,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m100001_0	),
Adb60111010101	(	adb60111010101,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m100001_0	),
Adb60111010110	(	adb60111010110,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m100001_0	),
Adb60111010111	(	adb60111010111,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m100001_0	),
Adb60111011000	(	adb60111011000,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m100001_0	),
Adb60111011001	(	adb60111011001,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m100001_0	),
Adb60111011010	(	adb60111011010,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m100001_0	),
Adb60111011011	(	adb60111011011,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m100001_0	),
Adb60111011100	(	adb60111011100,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m100001_0	),
Adb60111011101	(	adb60111011101,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m100001_0	),
Adb60111011110	(	adb60111011110,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m100001_0	),
Adb60111011111	(	adb60111011111,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m100001_0	),
Adb60111100000	(	adb60111100000,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m100001_0	),
Adb60111100001	(	adb60111100001,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m100001_0	),
Adb60111100010	(	adb60111100010,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m100001_0	),
Adb60111100011	(	adb60111100011,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m100001_0	),
Adb60111100100	(	adb60111100100,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m100001_0	),
Adb60111100101	(	adb60111100101,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m100001_0	),
Adb60111100110	(	adb60111100110,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m100001_0	),
Adb60111100111	(	adb60111100111,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m100001_0	),
Adb60111101000	(	adb60111101000,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m100001_0	),
Adb60111101001	(	adb60111101001,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m100001_0	),
Adb60111101010	(	adb60111101010,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m100001_0	),
Adb60111101011	(	adb60111101011,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m100001_0	),
Adb60111101100	(	adb60111101100,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m100001_0	),
Adb60111101101	(	adb60111101101,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m100001_0	),
Adb60111101110	(	adb60111101110,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m100001_0	),
Adb60111101111	(	adb60111101111,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m100001_0	),
Adb60111110000	(	adb60111110000,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m100001_0	),
Adb60111110001	(	adb60111110001,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m100001_0	),
Adb60111110010	(	adb60111110010,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m100001_0	),
Adb60111110011	(	adb60111110011,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m100001_0	),
Adb60111110100	(	adb60111110100,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m100001_0	),
Adb60111110101	(	adb60111110101,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m100001_0	),
Adb60111110110	(	adb60111110110,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m100001_0	),
Adb60111110111	(	adb60111110111,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m100001_0	),
Adb60111111000	(	adb60111111000,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m100001_0	),
Adb60111111001	(	adb60111111001,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m100001_0	),
Adb60111111010	(	adb60111111010,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m100001_0	),
Adb60111111011	(	adb60111111011,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m100001_0	),
Adb60111111100	(	adb60111111100,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m100001_0	),
Adb60111111101	(	adb60111111101,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m100001_0	),
Adb60111111110	(	adb60111111110,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m100001_0	),
Adb60111111111	(	adb60111111111,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m100001_0	),
Adb61000000000	(	adb61000000000,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m011001_0	),
Adb61000000001	(	adb61000000001,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m011001_0	),
Adb61000000010	(	adb61000000010,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m011001_0	),
Adb61000000011	(	adb61000000011,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m011001_0	),
Adb61000000100	(	adb61000000100,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m011001_0	),
Adb61000000101	(	adb61000000101,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m011001_0	),
Adb61000000110	(	adb61000000110,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m011001_0	),
Adb61000000111	(	adb61000000111,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m011001_0	),
Adb61000001000	(	adb61000001000,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m011001_0	),
Adb61000001001	(	adb61000001001,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m011001_0	),
Adb61000001010	(	adb61000001010,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m011001_0	),
Adb61000001011	(	adb61000001011,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m011001_0	),
Adb61000001100	(	adb61000001100,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m011001_0	),
Adb61000001101	(	adb61000001101,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m011001_0	),
Adb61000001110	(	adb61000001110,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m011001_0	),
Adb61000001111	(	adb61000001111,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m011001_0	),
Adb61000010000	(	adb61000010000,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m011001_0	),
Adb61000010001	(	adb61000010001,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m011001_0	),
Adb61000010010	(	adb61000010010,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m011001_0	),
Adb61000010011	(	adb61000010011,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m011001_0	),
Adb61000010100	(	adb61000010100,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m011001_0	),
Adb61000010101	(	adb61000010101,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m011001_0	),
Adb61000010110	(	adb61000010110,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m011001_0	),
Adb61000010111	(	adb61000010111,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m011001_0	),
Adb61000011000	(	adb61000011000,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m011001_0	),
Adb61000011001	(	adb61000011001,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m011001_0	),
Adb61000011010	(	adb61000011010,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m011001_0	),
Adb61000011011	(	adb61000011011,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m011001_0	),
Adb61000011100	(	adb61000011100,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m011001_0	),
Adb61000011101	(	adb61000011101,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m011001_0	),
Adb61000011110	(	adb61000011110,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m011001_0	),
Adb61000011111	(	adb61000011111,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m011001_0	),
Adb61000100000	(	adb61000100000,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m011001_0	),
Adb61000100001	(	adb61000100001,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m011001_0	),
Adb61000100010	(	adb61000100010,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m011001_0	),
Adb61000100011	(	adb61000100011,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m011001_0	),
Adb61000100100	(	adb61000100100,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m011001_0	),
Adb61000100101	(	adb61000100101,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m011001_0	),
Adb61000100110	(	adb61000100110,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m011001_0	),
Adb61000100111	(	adb61000100111,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m011001_0	),
Adb61000101000	(	adb61000101000,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m011001_0	),
Adb61000101001	(	adb61000101001,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m011001_0	),
Adb61000101010	(	adb61000101010,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m011001_0	),
Adb61000101011	(	adb61000101011,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m011001_0	),
Adb61000101100	(	adb61000101100,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m011001_0	),
Adb61000101101	(	adb61000101101,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m011001_0	),
Adb61000101110	(	adb61000101110,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m011001_0	),
Adb61000101111	(	adb61000101111,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m011001_0	),
Adb61000110000	(	adb61000110000,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m011001_0	),
Adb61000110001	(	adb61000110001,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m011001_0	),
Adb61000110010	(	adb61000110010,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m011001_0	),
Adb61000110011	(	adb61000110011,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m011001_0	),
Adb61000110100	(	adb61000110100,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m011001_0	),
Adb61000110101	(	adb61000110101,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m011001_0	),
Adb61000110110	(	adb61000110110,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m011001_0	),
Adb61000110111	(	adb61000110111,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m011001_0	),
Adb61000111000	(	adb61000111000,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m011001_0	),
Adb61000111001	(	adb61000111001,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m011001_0	),
Adb61000111010	(	adb61000111010,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m011001_0	),
Adb61000111011	(	adb61000111011,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m011001_0	),
Adb61000111100	(	adb61000111100,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m011001_0	),
Adb61000111101	(	adb61000111101,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m011001_0	),
Adb61000111110	(	adb61000111110,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m011001_0	),
Adb61000111111	(	adb61000111111,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m011001_0	),
Adb61001000000	(	adb61001000000,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m011001_0	),
Adb61001000001	(	adb61001000001,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m011001_0	),
Adb61001000010	(	adb61001000010,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m011001_0	),
Adb61001000011	(	adb61001000011,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m011001_0	),
Adb61001000100	(	adb61001000100,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m011001_0	),
Adb61001000101	(	adb61001000101,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m011001_0	),
Adb61001000110	(	adb61001000110,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m011001_0	),
Adb61001000111	(	adb61001000111,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m011001_0	),
Adb61001001000	(	adb61001001000,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m011001_0	),
Adb61001001001	(	adb61001001001,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m011001_0	),
Adb61001001010	(	adb61001001010,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m011001_0	),
Adb61001001011	(	adb61001001011,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m011001_0	),
Adb61001001100	(	adb61001001100,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m011001_0	),
Adb61001001101	(	adb61001001101,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m011001_0	),
Adb61001001110	(	adb61001001110,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m011001_0	),
Adb61001001111	(	adb61001001111,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m011001_0	),
Adb61001010000	(	adb61001010000,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m011001_0	),
Adb61001010001	(	adb61001010001,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m011001_0	),
Adb61001010010	(	adb61001010010,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m011001_0	),
Adb61001010011	(	adb61001010011,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m011001_0	),
Adb61001010100	(	adb61001010100,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m011001_0	),
Adb61001010101	(	adb61001010101,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m011001_0	),
Adb61001010110	(	adb61001010110,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m011001_0	),
Adb61001010111	(	adb61001010111,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m011001_0	),
Adb61001011000	(	adb61001011000,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m011001_0	),
Adb61001011001	(	adb61001011001,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m011001_0	),
Adb61001011010	(	adb61001011010,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m011001_0	),
Adb61001011011	(	adb61001011011,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m011001_0	),
Adb61001011100	(	adb61001011100,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m011001_0	),
Adb61001011101	(	adb61001011101,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m011001_0	),
Adb61001011110	(	adb61001011110,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m011001_0	),
Adb61001011111	(	adb61001011111,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m011001_0	),
Adb61001100000	(	adb61001100000,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m011001_0	),
Adb61001100001	(	adb61001100001,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m011001_0	),
Adb61001100010	(	adb61001100010,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m011001_0	),
Adb61001100011	(	adb61001100011,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m011001_0	),
Adb61001100100	(	adb61001100100,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m011001_0	),
Adb61001100101	(	adb61001100101,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m011001_0	),
Adb61001100110	(	adb61001100110,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m011001_0	),
Adb61001100111	(	adb61001100111,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m011001_0	),
Adb61001101000	(	adb61001101000,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m011001_0	),
Adb61001101001	(	adb61001101001,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m011001_0	),
Adb61001101010	(	adb61001101010,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m011001_0	),
Adb61001101011	(	adb61001101011,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m011001_0	),
Adb61001101100	(	adb61001101100,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m011001_0	),
Adb61001101101	(	adb61001101101,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m011001_0	),
Adb61001101110	(	adb61001101110,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m011001_0	),
Adb61001101111	(	adb61001101111,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m011001_0	),
Adb61001110000	(	adb61001110000,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m011001_0	),
Adb61001110001	(	adb61001110001,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m011001_0	),
Adb61001110010	(	adb61001110010,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m011001_0	),
Adb61001110011	(	adb61001110011,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m011001_0	),
Adb61001110100	(	adb61001110100,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m011001_0	),
Adb61001110101	(	adb61001110101,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m011001_0	),
Adb61001110110	(	adb61001110110,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m011001_0	),
Adb61001110111	(	adb61001110111,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m011001_0	),
Adb61001111000	(	adb61001111000,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m011001_0	),
Adb61001111001	(	adb61001111001,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m011001_0	),
Adb61001111010	(	adb61001111010,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m011001_0	),
Adb61001111011	(	adb61001111011,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m011001_0	),
Adb61001111100	(	adb61001111100,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m011001_0	),
Adb61001111101	(	adb61001111101,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m011001_0	),
Adb61001111110	(	adb61001111110,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m011001_0	),
Adb61001111111	(	adb61001111111,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m011001_0	),
Adb61010000000	(	adb61010000000,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m010001_0	),
Adb61010000001	(	adb61010000001,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m010001_0	),
Adb61010000010	(	adb61010000010,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m010001_0	),
Adb61010000011	(	adb61010000011,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m010001_0	),
Adb61010000100	(	adb61010000100,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m010001_0	),
Adb61010000101	(	adb61010000101,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m010001_0	),
Adb61010000110	(	adb61010000110,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m010001_0	),
Adb61010000111	(	adb61010000111,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m010001_0	),
Adb61010001000	(	adb61010001000,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m010001_0	),
Adb61010001001	(	adb61010001001,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m010001_0	),
Adb61010001010	(	adb61010001010,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m010001_0	),
Adb61010001011	(	adb61010001011,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m010001_0	),
Adb61010001100	(	adb61010001100,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m010001_0	),
Adb61010001101	(	adb61010001101,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m010001_0	),
Adb61010001110	(	adb61010001110,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m010001_0	),
Adb61010001111	(	adb61010001111,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m010001_0	),
Adb61010010000	(	adb61010010000,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m010001_0	),
Adb61010010001	(	adb61010010001,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m010001_0	),
Adb61010010010	(	adb61010010010,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m010001_0	),
Adb61010010011	(	adb61010010011,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m010001_0	),
Adb61010010100	(	adb61010010100,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m010001_0	),
Adb61010010101	(	adb61010010101,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m010001_0	),
Adb61010010110	(	adb61010010110,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m010001_0	),
Adb61010010111	(	adb61010010111,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m010001_0	),
Adb61010011000	(	adb61010011000,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m010001_0	),
Adb61010011001	(	adb61010011001,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m010001_0	),
Adb61010011010	(	adb61010011010,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m010001_0	),
Adb61010011011	(	adb61010011011,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m010001_0	),
Adb61010011100	(	adb61010011100,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m010001_0	),
Adb61010011101	(	adb61010011101,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m010001_0	),
Adb61010011110	(	adb61010011110,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m010001_0	),
Adb61010011111	(	adb61010011111,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m010001_0	),
Adb61010100000	(	adb61010100000,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m010001_0	),
Adb61010100001	(	adb61010100001,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m010001_0	),
Adb61010100010	(	adb61010100010,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m010001_0	),
Adb61010100011	(	adb61010100011,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m010001_0	),
Adb61010100100	(	adb61010100100,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m010001_0	),
Adb61010100101	(	adb61010100101,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m010001_0	),
Adb61010100110	(	adb61010100110,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m010001_0	),
Adb61010100111	(	adb61010100111,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m010001_0	),
Adb61010101000	(	adb61010101000,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m010001_0	),
Adb61010101001	(	adb61010101001,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m010001_0	),
Adb61010101010	(	adb61010101010,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m010001_0	),
Adb61010101011	(	adb61010101011,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m010001_0	),
Adb61010101100	(	adb61010101100,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m010001_0	),
Adb61010101101	(	adb61010101101,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m010001_0	),
Adb61010101110	(	adb61010101110,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m010001_0	),
Adb61010101111	(	adb61010101111,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m010001_0	),
Adb61010110000	(	adb61010110000,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m010001_0	),
Adb61010110001	(	adb61010110001,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m010001_0	),
Adb61010110010	(	adb61010110010,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m010001_0	),
Adb61010110011	(	adb61010110011,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m010001_0	),
Adb61010110100	(	adb61010110100,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m010001_0	),
Adb61010110101	(	adb61010110101,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m010001_0	),
Adb61010110110	(	adb61010110110,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m010001_0	),
Adb61010110111	(	adb61010110111,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m010001_0	),
Adb61010111000	(	adb61010111000,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m010001_0	),
Adb61010111001	(	adb61010111001,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m010001_0	),
Adb61010111010	(	adb61010111010,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m010001_0	),
Adb61010111011	(	adb61010111011,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m010001_0	),
Adb61010111100	(	adb61010111100,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m010001_0	),
Adb61010111101	(	adb61010111101,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m010001_0	),
Adb61010111110	(	adb61010111110,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m010001_0	),
Adb61010111111	(	adb61010111111,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m010001_0	),
Adb61011000000	(	adb61011000000,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m010001_0	),
Adb61011000001	(	adb61011000001,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m010001_0	),
Adb61011000010	(	adb61011000010,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m010001_0	),
Adb61011000011	(	adb61011000011,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m010001_0	),
Adb61011000100	(	adb61011000100,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m010001_0	),
Adb61011000101	(	adb61011000101,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m010001_0	),
Adb61011000110	(	adb61011000110,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m010001_0	),
Adb61011000111	(	adb61011000111,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m010001_0	),
Adb61011001000	(	adb61011001000,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m010001_0	),
Adb61011001001	(	adb61011001001,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m010001_0	),
Adb61011001010	(	adb61011001010,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m010001_0	),
Adb61011001011	(	adb61011001011,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m010001_0	),
Adb61011001100	(	adb61011001100,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m010001_0	),
Adb61011001101	(	adb61011001101,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m010001_0	),
Adb61011001110	(	adb61011001110,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m010001_0	),
Adb61011001111	(	adb61011001111,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m010001_0	),
Adb61011010000	(	adb61011010000,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m010001_0	),
Adb61011010001	(	adb61011010001,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m010001_0	),
Adb61011010010	(	adb61011010010,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m010001_0	),
Adb61011010011	(	adb61011010011,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m010001_0	),
Adb61011010100	(	adb61011010100,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m010001_0	),
Adb61011010101	(	adb61011010101,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m010001_0	),
Adb61011010110	(	adb61011010110,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m010001_0	),
Adb61011010111	(	adb61011010111,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m010001_0	),
Adb61011011000	(	adb61011011000,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m010001_0	),
Adb61011011001	(	adb61011011001,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m010001_0	),
Adb61011011010	(	adb61011011010,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m010001_0	),
Adb61011011011	(	adb61011011011,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m010001_0	),
Adb61011011100	(	adb61011011100,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m010001_0	),
Adb61011011101	(	adb61011011101,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m010001_0	),
Adb61011011110	(	adb61011011110,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m010001_0	),
Adb61011011111	(	adb61011011111,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m010001_0	),
Adb61011100000	(	adb61011100000,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m010001_0	),
Adb61011100001	(	adb61011100001,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m010001_0	),
Adb61011100010	(	adb61011100010,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m010001_0	),
Adb61011100011	(	adb61011100011,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m010001_0	),
Adb61011100100	(	adb61011100100,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m010001_0	),
Adb61011100101	(	adb61011100101,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m010001_0	),
Adb61011100110	(	adb61011100110,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m010001_0	),
Adb61011100111	(	adb61011100111,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m010001_0	),
Adb61011101000	(	adb61011101000,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m010001_0	),
Adb61011101001	(	adb61011101001,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m010001_0	),
Adb61011101010	(	adb61011101010,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m010001_0	),
Adb61011101011	(	adb61011101011,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m010001_0	),
Adb61011101100	(	adb61011101100,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m010001_0	),
Adb61011101101	(	adb61011101101,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m010001_0	),
Adb61011101110	(	adb61011101110,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m010001_0	),
Adb61011101111	(	adb61011101111,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m010001_0	),
Adb61011110000	(	adb61011110000,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m010001_0	),
Adb61011110001	(	adb61011110001,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m010001_0	),
Adb61011110010	(	adb61011110010,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m010001_0	),
Adb61011110011	(	adb61011110011,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m010001_0	),
Adb61011110100	(	adb61011110100,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m010001_0	),
Adb61011110101	(	adb61011110101,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m010001_0	),
Adb61011110110	(	adb61011110110,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m010001_0	),
Adb61011110111	(	adb61011110111,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m010001_0	),
Adb61011111000	(	adb61011111000,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m010001_0	),
Adb61011111001	(	adb61011111001,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m010001_0	),
Adb61011111010	(	adb61011111010,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m010001_0	),
Adb61011111011	(	adb61011111011,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m010001_0	),
Adb61011111100	(	adb61011111100,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m010001_0	),
Adb61011111101	(	adb61011111101,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m010001_0	),
Adb61011111110	(	adb61011111110,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m010001_0	),
Adb61011111111	(	adb61011111111,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m010001_0	),
Adb61100000000	(	adb61100000000,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m001001_0	),
Adb61100000001	(	adb61100000001,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m001001_0	),
Adb61100000010	(	adb61100000010,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m001001_0	),
Adb61100000011	(	adb61100000011,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m001001_0	),
Adb61100000100	(	adb61100000100,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m001001_0	),
Adb61100000101	(	adb61100000101,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m001001_0	),
Adb61100000110	(	adb61100000110,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m001001_0	),
Adb61100000111	(	adb61100000111,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m001001_0	),
Adb61100001000	(	adb61100001000,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m001001_0	),
Adb61100001001	(	adb61100001001,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m001001_0	),
Adb61100001010	(	adb61100001010,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m001001_0	),
Adb61100001011	(	adb61100001011,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m001001_0	),
Adb61100001100	(	adb61100001100,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m001001_0	),
Adb61100001101	(	adb61100001101,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m001001_0	),
Adb61100001110	(	adb61100001110,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m001001_0	),
Adb61100001111	(	adb61100001111,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m001001_0	),
Adb61100010000	(	adb61100010000,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m001001_0	),
Adb61100010001	(	adb61100010001,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m001001_0	),
Adb61100010010	(	adb61100010010,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m001001_0	),
Adb61100010011	(	adb61100010011,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m001001_0	),
Adb61100010100	(	adb61100010100,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m001001_0	),
Adb61100010101	(	adb61100010101,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m001001_0	),
Adb61100010110	(	adb61100010110,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m001001_0	),
Adb61100010111	(	adb61100010111,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m001001_0	),
Adb61100011000	(	adb61100011000,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m001001_0	),
Adb61100011001	(	adb61100011001,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m001001_0	),
Adb61100011010	(	adb61100011010,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m001001_0	),
Adb61100011011	(	adb61100011011,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m001001_0	),
Adb61100011100	(	adb61100011100,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m001001_0	),
Adb61100011101	(	adb61100011101,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m001001_0	),
Adb61100011110	(	adb61100011110,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m001001_0	),
Adb61100011111	(	adb61100011111,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m001001_0	),
Adb61100100000	(	adb61100100000,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m001001_0	),
Adb61100100001	(	adb61100100001,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m001001_0	),
Adb61100100010	(	adb61100100010,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m001001_0	),
Adb61100100011	(	adb61100100011,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m001001_0	),
Adb61100100100	(	adb61100100100,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m001001_0	),
Adb61100100101	(	adb61100100101,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m001001_0	),
Adb61100100110	(	adb61100100110,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m001001_0	),
Adb61100100111	(	adb61100100111,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m001001_0	),
Adb61100101000	(	adb61100101000,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m001001_0	),
Adb61100101001	(	adb61100101001,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m001001_0	),
Adb61100101010	(	adb61100101010,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m001001_0	),
Adb61100101011	(	adb61100101011,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m001001_0	),
Adb61100101100	(	adb61100101100,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m001001_0	),
Adb61100101101	(	adb61100101101,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m001001_0	),
Adb61100101110	(	adb61100101110,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m001001_0	),
Adb61100101111	(	adb61100101111,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m001001_0	),
Adb61100110000	(	adb61100110000,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m001001_0	),
Adb61100110001	(	adb61100110001,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m001001_0	),
Adb61100110010	(	adb61100110010,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m001001_0	),
Adb61100110011	(	adb61100110011,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m001001_0	),
Adb61100110100	(	adb61100110100,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m001001_0	),
Adb61100110101	(	adb61100110101,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m001001_0	),
Adb61100110110	(	adb61100110110,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m001001_0	),
Adb61100110111	(	adb61100110111,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m001001_0	),
Adb61100111000	(	adb61100111000,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m001001_0	),
Adb61100111001	(	adb61100111001,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m001001_0	),
Adb61100111010	(	adb61100111010,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m001001_0	),
Adb61100111011	(	adb61100111011,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m001001_0	),
Adb61100111100	(	adb61100111100,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m001001_0	),
Adb61100111101	(	adb61100111101,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m001001_0	),
Adb61100111110	(	adb61100111110,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m001001_0	),
Adb61100111111	(	adb61100111111,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m001001_0	),
Adb61101000000	(	adb61101000000,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m001001_0	),
Adb61101000001	(	adb61101000001,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m001001_0	),
Adb61101000010	(	adb61101000010,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m001001_0	),
Adb61101000011	(	adb61101000011,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m001001_0	),
Adb61101000100	(	adb61101000100,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m001001_0	),
Adb61101000101	(	adb61101000101,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m001001_0	),
Adb61101000110	(	adb61101000110,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m001001_0	),
Adb61101000111	(	adb61101000111,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m001001_0	),
Adb61101001000	(	adb61101001000,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m001001_0	),
Adb61101001001	(	adb61101001001,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m001001_0	),
Adb61101001010	(	adb61101001010,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m001001_0	),
Adb61101001011	(	adb61101001011,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m001001_0	),
Adb61101001100	(	adb61101001100,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m001001_0	),
Adb61101001101	(	adb61101001101,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m001001_0	),
Adb61101001110	(	adb61101001110,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m001001_0	),
Adb61101001111	(	adb61101001111,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m001001_0	),
Adb61101010000	(	adb61101010000,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m001001_0	),
Adb61101010001	(	adb61101010001,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m001001_0	),
Adb61101010010	(	adb61101010010,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m001001_0	),
Adb61101010011	(	adb61101010011,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m001001_0	),
Adb61101010100	(	adb61101010100,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m001001_0	),
Adb61101010101	(	adb61101010101,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m001001_0	),
Adb61101010110	(	adb61101010110,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m001001_0	),
Adb61101010111	(	adb61101010111,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m001001_0	),
Adb61101011000	(	adb61101011000,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m001001_0	),
Adb61101011001	(	adb61101011001,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m001001_0	),
Adb61101011010	(	adb61101011010,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m001001_0	),
Adb61101011011	(	adb61101011011,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m001001_0	),
Adb61101011100	(	adb61101011100,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m001001_0	),
Adb61101011101	(	adb61101011101,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m001001_0	),
Adb61101011110	(	adb61101011110,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m001001_0	),
Adb61101011111	(	adb61101011111,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m001001_0	),
Adb61101100000	(	adb61101100000,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m001001_0	),
Adb61101100001	(	adb61101100001,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m001001_0	),
Adb61101100010	(	adb61101100010,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m001001_0	),
Adb61101100011	(	adb61101100011,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m001001_0	),
Adb61101100100	(	adb61101100100,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m001001_0	),
Adb61101100101	(	adb61101100101,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m001001_0	),
Adb61101100110	(	adb61101100110,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m001001_0	),
Adb61101100111	(	adb61101100111,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m001001_0	),
Adb61101101000	(	adb61101101000,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m001001_0	),
Adb61101101001	(	adb61101101001,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m001001_0	),
Adb61101101010	(	adb61101101010,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m001001_0	),
Adb61101101011	(	adb61101101011,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m001001_0	),
Adb61101101100	(	adb61101101100,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m001001_0	),
Adb61101101101	(	adb61101101101,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m001001_0	),
Adb61101101110	(	adb61101101110,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m001001_0	),
Adb61101101111	(	adb61101101111,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m001001_0	),
Adb61101110000	(	adb61101110000,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m001001_0	),
Adb61101110001	(	adb61101110001,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m001001_0	),
Adb61101110010	(	adb61101110010,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m001001_0	),
Adb61101110011	(	adb61101110011,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m001001_0	),
Adb61101110100	(	adb61101110100,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m001001_0	),
Adb61101110101	(	adb61101110101,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m001001_0	),
Adb61101110110	(	adb61101110110,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m001001_0	),
Adb61101110111	(	adb61101110111,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m001001_0	),
Adb61101111000	(	adb61101111000,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m001001_0	),
Adb61101111001	(	adb61101111001,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m001001_0	),
Adb61101111010	(	adb61101111010,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m001001_0	),
Adb61101111011	(	adb61101111011,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m001001_0	),
Adb61101111100	(	adb61101111100,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m001001_0	),
Adb61101111101	(	adb61101111101,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m001001_0	),
Adb61101111110	(	adb61101111110,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m001001_0	),
Adb61101111111	(	adb61101111111,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m001001_0	),
Adb61110000000	(	adb61110000000,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m000001_0	),
Adb61110000001	(	adb61110000001,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m000001_0	),
Adb61110000010	(	adb61110000010,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m000001_0	),
Adb61110000011	(	adb61110000011,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m000001_0	),
Adb61110000100	(	adb61110000100,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m000001_0	),
Adb61110000101	(	adb61110000101,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m000001_0	),
Adb61110000110	(	adb61110000110,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m000001_0	),
Adb61110000111	(	adb61110000111,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m000001_0	),
Adb61110001000	(	adb61110001000,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m000001_0	),
Adb61110001001	(	adb61110001001,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m000001_0	),
Adb61110001010	(	adb61110001010,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m000001_0	),
Adb61110001011	(	adb61110001011,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m000001_0	),
Adb61110001100	(	adb61110001100,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m000001_0	),
Adb61110001101	(	adb61110001101,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m000001_0	),
Adb61110001110	(	adb61110001110,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m000001_0	),
Adb61110001111	(	adb61110001111,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m000001_0	),
Adb61110010000	(	adb61110010000,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m000001_0	),
Adb61110010001	(	adb61110010001,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m000001_0	),
Adb61110010010	(	adb61110010010,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m000001_0	),
Adb61110010011	(	adb61110010011,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m000001_0	),
Adb61110010100	(	adb61110010100,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m000001_0	),
Adb61110010101	(	adb61110010101,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m000001_0	),
Adb61110010110	(	adb61110010110,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m000001_0	),
Adb61110010111	(	adb61110010111,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m000001_0	),
Adb61110011000	(	adb61110011000,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m000001_0	),
Adb61110011001	(	adb61110011001,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m000001_0	),
Adb61110011010	(	adb61110011010,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m000001_0	),
Adb61110011011	(	adb61110011011,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m000001_0	),
Adb61110011100	(	adb61110011100,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m000001_0	),
Adb61110011101	(	adb61110011101,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m000001_0	),
Adb61110011110	(	adb61110011110,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m000001_0	),
Adb61110011111	(	adb61110011111,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m000001_0	),
Adb61110100000	(	adb61110100000,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m000001_0	),
Adb61110100001	(	adb61110100001,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m000001_0	),
Adb61110100010	(	adb61110100010,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m000001_0	),
Adb61110100011	(	adb61110100011,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m000001_0	),
Adb61110100100	(	adb61110100100,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m000001_0	),
Adb61110100101	(	adb61110100101,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m000001_0	),
Adb61110100110	(	adb61110100110,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m000001_0	),
Adb61110100111	(	adb61110100111,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m000001_0	),
Adb61110101000	(	adb61110101000,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m000001_0	),
Adb61110101001	(	adb61110101001,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m000001_0	),
Adb61110101010	(	adb61110101010,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m000001_0	),
Adb61110101011	(	adb61110101011,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m000001_0	),
Adb61110101100	(	adb61110101100,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m000001_0	),
Adb61110101101	(	adb61110101101,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m000001_0	),
Adb61110101110	(	adb61110101110,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m000001_0	),
Adb61110101111	(	adb61110101111,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m000001_0	),
Adb61110110000	(	adb61110110000,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m000001_0	),
Adb61110110001	(	adb61110110001,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m000001_0	),
Adb61110110010	(	adb61110110010,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m000001_0	),
Adb61110110011	(	adb61110110011,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m000001_0	),
Adb61110110100	(	adb61110110100,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m000001_0	),
Adb61110110101	(	adb61110110101,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m000001_0	),
Adb61110110110	(	adb61110110110,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m000001_0	),
Adb61110110111	(	adb61110110111,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m000001_0	),
Adb61110111000	(	adb61110111000,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m000001_0	),
Adb61110111001	(	adb61110111001,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m000001_0	),
Adb61110111010	(	adb61110111010,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m000001_0	),
Adb61110111011	(	adb61110111011,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m000001_0	),
Adb61110111100	(	adb61110111100,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m000001_0	),
Adb61110111101	(	adb61110111101,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m000001_0	),
Adb61110111110	(	adb61110111110,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m000001_0	),
Adb61110111111	(	adb61110111111,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m000001_0	),
Adb61111000000	(	adb61111000000,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m000001_0	),
Adb61111000001	(	adb61111000001,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m000001_0	),
Adb61111000010	(	adb61111000010,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m000001_0	),
Adb61111000011	(	adb61111000011,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m000001_0	),
Adb61111000100	(	adb61111000100,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m000001_0	),
Adb61111000101	(	adb61111000101,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m000001_0	),
Adb61111000110	(	adb61111000110,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m000001_0	),
Adb61111000111	(	adb61111000111,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m000001_0	),
Adb61111001000	(	adb61111001000,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m000001_0	),
Adb61111001001	(	adb61111001001,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m000001_0	),
Adb61111001010	(	adb61111001010,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m000001_0	),
Adb61111001011	(	adb61111001011,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m000001_0	),
Adb61111001100	(	adb61111001100,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m000001_0	),
Adb61111001101	(	adb61111001101,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m000001_0	),
Adb61111001110	(	adb61111001110,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m000001_0	),
Adb61111001111	(	adb61111001111,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m000001_0	),
Adb61111010000	(	adb61111010000,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m000001_0	),
Adb61111010001	(	adb61111010001,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m000001_0	),
Adb61111010010	(	adb61111010010,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m000001_0	),
Adb61111010011	(	adb61111010011,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m000001_0	),
Adb61111010100	(	adb61111010100,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m000001_0	),
Adb61111010101	(	adb61111010101,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m000001_0	),
Adb61111010110	(	adb61111010110,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m000001_0	),
Adb61111010111	(	adb61111010111,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m000001_0	),
Adb61111011000	(	adb61111011000,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m000001_0	),
Adb61111011001	(	adb61111011001,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m000001_0	),
Adb61111011010	(	adb61111011010,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m000001_0	),
Adb61111011011	(	adb61111011011,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m000001_0	),
Adb61111011100	(	adb61111011100,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m000001_0	),
Adb61111011101	(	adb61111011101,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m000001_0	),
Adb61111011110	(	adb61111011110,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m000001_0	),
Adb61111011111	(	adb61111011111,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m000001_0	),
Adb61111100000	(	adb61111100000,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m000001_0	),
Adb61111100001	(	adb61111100001,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m000001_0	),
Adb61111100010	(	adb61111100010,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m000001_0	),
Adb61111100011	(	adb61111100011,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m000001_0	),
Adb61111100100	(	adb61111100100,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m000001_0	),
Adb61111100101	(	adb61111100101,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m000001_0	),
Adb61111100110	(	adb61111100110,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m000001_0	),
Adb61111100111	(	adb61111100111,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m000001_0	),
Adb61111101000	(	adb61111101000,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m000001_0	),
Adb61111101001	(	adb61111101001,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m000001_0	),
Adb61111101010	(	adb61111101010,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m000001_0	),
Adb61111101011	(	adb61111101011,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m000001_0	),
Adb61111101100	(	adb61111101100,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m000001_0	),
Adb61111101101	(	adb61111101101,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m000001_0	),
Adb61111101110	(	adb61111101110,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m000001_0	),
Adb61111101111	(	adb61111101111,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m000001_0	),
Adb61111110000	(	adb61111110000,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m000001_0	),
Adb61111110001	(	adb61111110001,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m000001_0	),
Adb61111110010	(	adb61111110010,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m000001_0	),
Adb61111110011	(	adb61111110011,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m000001_0	),
Adb61111110100	(	adb61111110100,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m000001_0	),
Adb61111110101	(	adb61111110101,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m000001_0	),
Adb61111110110	(	adb61111110110,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m000001_0	),
Adb61111110111	(	adb61111110111,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m000001_0	),
Adb61111111000	(	adb61111111000,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m000001_0	),
Adb61111111001	(	adb61111111001,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m000001_0	),
Adb61111111010	(	adb61111111010,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m000001_0	),
Adb61111111011	(	adb61111111011,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m000001_0	),
Adb61111111100	(	adb61111111100,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m000001_0	),
Adb61111111101	(	adb61111111101,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m000001_0	),
Adb61111111110	(	adb61111111110,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m000001_0	),
Adb61111111111	(	adb61111111111,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m000001_0	),
       Adb700(adb700,n0011,n0010,n0009,m0010),
       Adb701(adb701,n0011,n0010,m0009,m0010),
       Adb710(adb710,n0011,m0010,n0009,m0010),
       Adb711(adb711,n0011,m0010,m0009,m0010),
Adb70000000000	(	adb70000000000,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m111000_0	),
Adb70000000001	(	adb70000000001,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m111000_0	),
Adb70000000010	(	adb70000000010,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m111000_0	),
Adb70000000011	(	adb70000000011,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m111000_0	),
Adb70000000100	(	adb70000000100,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m111000_0	),
Adb70000000101	(	adb70000000101,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m111000_0	),
Adb70000000110	(	adb70000000110,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m111000_0	),
Adb70000000111	(	adb70000000111,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m111000_0	),
Adb70000001000	(	adb70000001000,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m111000_0	),
Adb70000001001	(	adb70000001001,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m111000_0	),
Adb70000001010	(	adb70000001010,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m111000_0	),
Adb70000001011	(	adb70000001011,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m111000_0	),
Adb70000001100	(	adb70000001100,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m111000_0	),
Adb70000001101	(	adb70000001101,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m111000_0	),
Adb70000001110	(	adb70000001110,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m111000_0	),
Adb70000001111	(	adb70000001111,	n0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m111000_0	),
Adb70000010000	(	adb70000010000,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m111000_0	),
Adb70000010001	(	adb70000010001,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m111000_0	),
Adb70000010010	(	adb70000010010,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m111000_0	),
Adb70000010011	(	adb70000010011,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m111000_0	),
Adb70000010100	(	adb70000010100,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m111000_0	),
Adb70000010101	(	adb70000010101,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m111000_0	),
Adb70000010110	(	adb70000010110,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m111000_0	),
Adb70000010111	(	adb70000010111,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m111000_0	),
Adb70000011000	(	adb70000011000,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m111000_0	),
Adb70000011001	(	adb70000011001,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m111000_0	),
Adb70000011010	(	adb70000011010,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m111000_0	),
Adb70000011011	(	adb70000011011,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m111000_0	),
Adb70000011100	(	adb70000011100,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m111000_0	),
Adb70000011101	(	adb70000011101,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m111000_0	),
Adb70000011110	(	adb70000011110,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m111000_0	),
Adb70000011111	(	adb70000011111,	n0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m111000_0	),
Adb70000100000	(	adb70000100000,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m111000_0	),
Adb70000100001	(	adb70000100001,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m111000_0	),
Adb70000100010	(	adb70000100010,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m111000_0	),
Adb70000100011	(	adb70000100011,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m111000_0	),
Adb70000100100	(	adb70000100100,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m111000_0	),
Adb70000100101	(	adb70000100101,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m111000_0	),
Adb70000100110	(	adb70000100110,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m111000_0	),
Adb70000100111	(	adb70000100111,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m111000_0	),
Adb70000101000	(	adb70000101000,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m111000_0	),
Adb70000101001	(	adb70000101001,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m111000_0	),
Adb70000101010	(	adb70000101010,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m111000_0	),
Adb70000101011	(	adb70000101011,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m111000_0	),
Adb70000101100	(	adb70000101100,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m111000_0	),
Adb70000101101	(	adb70000101101,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m111000_0	),
Adb70000101110	(	adb70000101110,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m111000_0	),
Adb70000101111	(	adb70000101111,	n0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m111000_0	),
Adb70000110000	(	adb70000110000,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m111000_0	),
Adb70000110001	(	adb70000110001,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m111000_0	),
Adb70000110010	(	adb70000110010,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m111000_0	),
Adb70000110011	(	adb70000110011,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m111000_0	),
Adb70000110100	(	adb70000110100,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m111000_0	),
Adb70000110101	(	adb70000110101,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m111000_0	),
Adb70000110110	(	adb70000110110,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m111000_0	),
Adb70000110111	(	adb70000110111,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m111000_0	),
Adb70000111000	(	adb70000111000,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m111000_0	),
Adb70000111001	(	adb70000111001,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m111000_0	),
Adb70000111010	(	adb70000111010,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m111000_0	),
Adb70000111011	(	adb70000111011,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m111000_0	),
Adb70000111100	(	adb70000111100,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m111000_0	),
Adb70000111101	(	adb70000111101,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m111000_0	),
Adb70000111110	(	adb70000111110,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m111000_0	),
Adb70000111111	(	adb70000111111,	n0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m111000_0	),
Adb70001000000	(	adb70001000000,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m111000_0	),
Adb70001000001	(	adb70001000001,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m111000_0	),
Adb70001000010	(	adb70001000010,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m111000_0	),
Adb70001000011	(	adb70001000011,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m111000_0	),
Adb70001000100	(	adb70001000100,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m111000_0	),
Adb70001000101	(	adb70001000101,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m111000_0	),
Adb70001000110	(	adb70001000110,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m111000_0	),
Adb70001000111	(	adb70001000111,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m111000_0	),
Adb70001001000	(	adb70001001000,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m111000_0	),
Adb70001001001	(	adb70001001001,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m111000_0	),
Adb70001001010	(	adb70001001010,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m111000_0	),
Adb70001001011	(	adb70001001011,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m111000_0	),
Adb70001001100	(	adb70001001100,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m111000_0	),
Adb70001001101	(	adb70001001101,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m111000_0	),
Adb70001001110	(	adb70001001110,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m111000_0	),
Adb70001001111	(	adb70001001111,	n0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m111000_0	),
Adb70001010000	(	adb70001010000,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m111000_0	),
Adb70001010001	(	adb70001010001,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m111000_0	),
Adb70001010010	(	adb70001010010,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m111000_0	),
Adb70001010011	(	adb70001010011,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m111000_0	),
Adb70001010100	(	adb70001010100,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m111000_0	),
Adb70001010101	(	adb70001010101,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m111000_0	),
Adb70001010110	(	adb70001010110,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m111000_0	),
Adb70001010111	(	adb70001010111,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m111000_0	),
Adb70001011000	(	adb70001011000,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m111000_0	),
Adb70001011001	(	adb70001011001,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m111000_0	),
Adb70001011010	(	adb70001011010,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m111000_0	),
Adb70001011011	(	adb70001011011,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m111000_0	),
Adb70001011100	(	adb70001011100,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m111000_0	),
Adb70001011101	(	adb70001011101,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m111000_0	),
Adb70001011110	(	adb70001011110,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m111000_0	),
Adb70001011111	(	adb70001011111,	n0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m111000_0	),
Adb70001100000	(	adb70001100000,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m111000_0	),
Adb70001100001	(	adb70001100001,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m111000_0	),
Adb70001100010	(	adb70001100010,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m111000_0	),
Adb70001100011	(	adb70001100011,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m111000_0	),
Adb70001100100	(	adb70001100100,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m111000_0	),
Adb70001100101	(	adb70001100101,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m111000_0	),
Adb70001100110	(	adb70001100110,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m111000_0	),
Adb70001100111	(	adb70001100111,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m111000_0	),
Adb70001101000	(	adb70001101000,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m111000_0	),
Adb70001101001	(	adb70001101001,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m111000_0	),
Adb70001101010	(	adb70001101010,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m111000_0	),
Adb70001101011	(	adb70001101011,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m111000_0	),
Adb70001101100	(	adb70001101100,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m111000_0	),
Adb70001101101	(	adb70001101101,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m111000_0	),
Adb70001101110	(	adb70001101110,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m111000_0	),
Adb70001101111	(	adb70001101111,	n0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m111000_0	),
Adb70001110000	(	adb70001110000,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m111000_0	),
Adb70001110001	(	adb70001110001,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m111000_0	),
Adb70001110010	(	adb70001110010,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m111000_0	),
Adb70001110011	(	adb70001110011,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m111000_0	),
Adb70001110100	(	adb70001110100,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m111000_0	),
Adb70001110101	(	adb70001110101,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m111000_0	),
Adb70001110110	(	adb70001110110,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m111000_0	),
Adb70001110111	(	adb70001110111,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m111000_0	),
Adb70001111000	(	adb70001111000,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m111000_0	),
Adb70001111001	(	adb70001111001,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m111000_0	),
Adb70001111010	(	adb70001111010,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m111000_0	),
Adb70001111011	(	adb70001111011,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m111000_0	),
Adb70001111100	(	adb70001111100,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m111000_0	),
Adb70001111101	(	adb70001111101,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m111000_0	),
Adb70001111110	(	adb70001111110,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m111000_0	),
Adb70001111111	(	adb70001111111,	n0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m111000_0	),
Adb70010000000	(	adb70010000000,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m110000_0	),
Adb70010000001	(	adb70010000001,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m110000_0	),
Adb70010000010	(	adb70010000010,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m110000_0	),
Adb70010000011	(	adb70010000011,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m110000_0	),
Adb70010000100	(	adb70010000100,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m110000_0	),
Adb70010000101	(	adb70010000101,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m110000_0	),
Adb70010000110	(	adb70010000110,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m110000_0	),
Adb70010000111	(	adb70010000111,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m110000_0	),
Adb70010001000	(	adb70010001000,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m110000_0	),
Adb70010001001	(	adb70010001001,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m110000_0	),
Adb70010001010	(	adb70010001010,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m110000_0	),
Adb70010001011	(	adb70010001011,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m110000_0	),
Adb70010001100	(	adb70010001100,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m110000_0	),
Adb70010001101	(	adb70010001101,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m110000_0	),
Adb70010001110	(	adb70010001110,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m110000_0	),
Adb70010001111	(	adb70010001111,	n0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m110000_0	),
Adb70010010000	(	adb70010010000,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m110000_0	),
Adb70010010001	(	adb70010010001,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m110000_0	),
Adb70010010010	(	adb70010010010,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m110000_0	),
Adb70010010011	(	adb70010010011,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m110000_0	),
Adb70010010100	(	adb70010010100,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m110000_0	),
Adb70010010101	(	adb70010010101,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m110000_0	),
Adb70010010110	(	adb70010010110,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m110000_0	),
Adb70010010111	(	adb70010010111,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m110000_0	),
Adb70010011000	(	adb70010011000,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m110000_0	),
Adb70010011001	(	adb70010011001,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m110000_0	),
Adb70010011010	(	adb70010011010,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m110000_0	),
Adb70010011011	(	adb70010011011,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m110000_0	),
Adb70010011100	(	adb70010011100,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m110000_0	),
Adb70010011101	(	adb70010011101,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m110000_0	),
Adb70010011110	(	adb70010011110,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m110000_0	),
Adb70010011111	(	adb70010011111,	n0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m110000_0	),
Adb70010100000	(	adb70010100000,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m110000_0	),
Adb70010100001	(	adb70010100001,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m110000_0	),
Adb70010100010	(	adb70010100010,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m110000_0	),
Adb70010100011	(	adb70010100011,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m110000_0	),
Adb70010100100	(	adb70010100100,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m110000_0	),
Adb70010100101	(	adb70010100101,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m110000_0	),
Adb70010100110	(	adb70010100110,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m110000_0	),
Adb70010100111	(	adb70010100111,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m110000_0	),
Adb70010101000	(	adb70010101000,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m110000_0	),
Adb70010101001	(	adb70010101001,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m110000_0	),
Adb70010101010	(	adb70010101010,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m110000_0	),
Adb70010101011	(	adb70010101011,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m110000_0	),
Adb70010101100	(	adb70010101100,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m110000_0	),
Adb70010101101	(	adb70010101101,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m110000_0	),
Adb70010101110	(	adb70010101110,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m110000_0	),
Adb70010101111	(	adb70010101111,	n0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m110000_0	),
Adb70010110000	(	adb70010110000,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m110000_0	),
Adb70010110001	(	adb70010110001,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m110000_0	),
Adb70010110010	(	adb70010110010,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m110000_0	),
Adb70010110011	(	adb70010110011,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m110000_0	),
Adb70010110100	(	adb70010110100,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m110000_0	),
Adb70010110101	(	adb70010110101,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m110000_0	),
Adb70010110110	(	adb70010110110,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m110000_0	),
Adb70010110111	(	adb70010110111,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m110000_0	),
Adb70010111000	(	adb70010111000,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m110000_0	),
Adb70010111001	(	adb70010111001,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m110000_0	),
Adb70010111010	(	adb70010111010,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m110000_0	),
Adb70010111011	(	adb70010111011,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m110000_0	),
Adb70010111100	(	adb70010111100,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m110000_0	),
Adb70010111101	(	adb70010111101,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m110000_0	),
Adb70010111110	(	adb70010111110,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m110000_0	),
Adb70010111111	(	adb70010111111,	n0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m110000_0	),
Adb70011000000	(	adb70011000000,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m110000_0	),
Adb70011000001	(	adb70011000001,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m110000_0	),
Adb70011000010	(	adb70011000010,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m110000_0	),
Adb70011000011	(	adb70011000011,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m110000_0	),
Adb70011000100	(	adb70011000100,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m110000_0	),
Adb70011000101	(	adb70011000101,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m110000_0	),
Adb70011000110	(	adb70011000110,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m110000_0	),
Adb70011000111	(	adb70011000111,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m110000_0	),
Adb70011001000	(	adb70011001000,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m110000_0	),
Adb70011001001	(	adb70011001001,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m110000_0	),
Adb70011001010	(	adb70011001010,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m110000_0	),
Adb70011001011	(	adb70011001011,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m110000_0	),
Adb70011001100	(	adb70011001100,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m110000_0	),
Adb70011001101	(	adb70011001101,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m110000_0	),
Adb70011001110	(	adb70011001110,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m110000_0	),
Adb70011001111	(	adb70011001111,	n0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m110000_0	),
Adb70011010000	(	adb70011010000,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m110000_0	),
Adb70011010001	(	adb70011010001,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m110000_0	),
Adb70011010010	(	adb70011010010,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m110000_0	),
Adb70011010011	(	adb70011010011,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m110000_0	),
Adb70011010100	(	adb70011010100,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m110000_0	),
Adb70011010101	(	adb70011010101,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m110000_0	),
Adb70011010110	(	adb70011010110,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m110000_0	),
Adb70011010111	(	adb70011010111,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m110000_0	),
Adb70011011000	(	adb70011011000,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m110000_0	),
Adb70011011001	(	adb70011011001,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m110000_0	),
Adb70011011010	(	adb70011011010,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m110000_0	),
Adb70011011011	(	adb70011011011,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m110000_0	),
Adb70011011100	(	adb70011011100,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m110000_0	),
Adb70011011101	(	adb70011011101,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m110000_0	),
Adb70011011110	(	adb70011011110,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m110000_0	),
Adb70011011111	(	adb70011011111,	n0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m110000_0	),
Adb70011100000	(	adb70011100000,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m110000_0	),
Adb70011100001	(	adb70011100001,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m110000_0	),
Adb70011100010	(	adb70011100010,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m110000_0	),
Adb70011100011	(	adb70011100011,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m110000_0	),
Adb70011100100	(	adb70011100100,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m110000_0	),
Adb70011100101	(	adb70011100101,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m110000_0	),
Adb70011100110	(	adb70011100110,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m110000_0	),
Adb70011100111	(	adb70011100111,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m110000_0	),
Adb70011101000	(	adb70011101000,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m110000_0	),
Adb70011101001	(	adb70011101001,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m110000_0	),
Adb70011101010	(	adb70011101010,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m110000_0	),
Adb70011101011	(	adb70011101011,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m110000_0	),
Adb70011101100	(	adb70011101100,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m110000_0	),
Adb70011101101	(	adb70011101101,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m110000_0	),
Adb70011101110	(	adb70011101110,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m110000_0	),
Adb70011101111	(	adb70011101111,	n0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m110000_0	),
Adb70011110000	(	adb70011110000,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m110000_0	),
Adb70011110001	(	adb70011110001,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m110000_0	),
Adb70011110010	(	adb70011110010,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m110000_0	),
Adb70011110011	(	adb70011110011,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m110000_0	),
Adb70011110100	(	adb70011110100,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m110000_0	),
Adb70011110101	(	adb70011110101,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m110000_0	),
Adb70011110110	(	adb70011110110,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m110000_0	),
Adb70011110111	(	adb70011110111,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m110000_0	),
Adb70011111000	(	adb70011111000,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m110000_0	),
Adb70011111001	(	adb70011111001,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m110000_0	),
Adb70011111010	(	adb70011111010,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m110000_0	),
Adb70011111011	(	adb70011111011,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m110000_0	),
Adb70011111100	(	adb70011111100,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m110000_0	),
Adb70011111101	(	adb70011111101,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m110000_0	),
Adb70011111110	(	adb70011111110,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m110000_0	),
Adb70011111111	(	adb70011111111,	n0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m110000_0	),
Adb70100000000	(	adb70100000000,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m101000_0	),
Adb70100000001	(	adb70100000001,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m101000_0	),
Adb70100000010	(	adb70100000010,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m101000_0	),
Adb70100000011	(	adb70100000011,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m101000_0	),
Adb70100000100	(	adb70100000100,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m101000_0	),
Adb70100000101	(	adb70100000101,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m101000_0	),
Adb70100000110	(	adb70100000110,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m101000_0	),
Adb70100000111	(	adb70100000111,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m101000_0	),
Adb70100001000	(	adb70100001000,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m101000_0	),
Adb70100001001	(	adb70100001001,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m101000_0	),
Adb70100001010	(	adb70100001010,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m101000_0	),
Adb70100001011	(	adb70100001011,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m101000_0	),
Adb70100001100	(	adb70100001100,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m101000_0	),
Adb70100001101	(	adb70100001101,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m101000_0	),
Adb70100001110	(	adb70100001110,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m101000_0	),
Adb70100001111	(	adb70100001111,	n0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m101000_0	),
Adb70100010000	(	adb70100010000,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m101000_0	),
Adb70100010001	(	adb70100010001,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m101000_0	),
Adb70100010010	(	adb70100010010,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m101000_0	),
Adb70100010011	(	adb70100010011,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m101000_0	),
Adb70100010100	(	adb70100010100,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m101000_0	),
Adb70100010101	(	adb70100010101,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m101000_0	),
Adb70100010110	(	adb70100010110,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m101000_0	),
Adb70100010111	(	adb70100010111,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m101000_0	),
Adb70100011000	(	adb70100011000,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m101000_0	),
Adb70100011001	(	adb70100011001,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m101000_0	),
Adb70100011010	(	adb70100011010,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m101000_0	),
Adb70100011011	(	adb70100011011,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m101000_0	),
Adb70100011100	(	adb70100011100,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m101000_0	),
Adb70100011101	(	adb70100011101,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m101000_0	),
Adb70100011110	(	adb70100011110,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m101000_0	),
Adb70100011111	(	adb70100011111,	n0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m101000_0	),
Adb70100100000	(	adb70100100000,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m101000_0	),
Adb70100100001	(	adb70100100001,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m101000_0	),
Adb70100100010	(	adb70100100010,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m101000_0	),
Adb70100100011	(	adb70100100011,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m101000_0	),
Adb70100100100	(	adb70100100100,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m101000_0	),
Adb70100100101	(	adb70100100101,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m101000_0	),
Adb70100100110	(	adb70100100110,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m101000_0	),
Adb70100100111	(	adb70100100111,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m101000_0	),
Adb70100101000	(	adb70100101000,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m101000_0	),
Adb70100101001	(	adb70100101001,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m101000_0	),
Adb70100101010	(	adb70100101010,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m101000_0	),
Adb70100101011	(	adb70100101011,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m101000_0	),
Adb70100101100	(	adb70100101100,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m101000_0	),
Adb70100101101	(	adb70100101101,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m101000_0	),
Adb70100101110	(	adb70100101110,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m101000_0	),
Adb70100101111	(	adb70100101111,	n0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m101000_0	),
Adb70100110000	(	adb70100110000,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m101000_0	),
Adb70100110001	(	adb70100110001,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m101000_0	),
Adb70100110010	(	adb70100110010,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m101000_0	),
Adb70100110011	(	adb70100110011,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m101000_0	),
Adb70100110100	(	adb70100110100,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m101000_0	),
Adb70100110101	(	adb70100110101,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m101000_0	),
Adb70100110110	(	adb70100110110,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m101000_0	),
Adb70100110111	(	adb70100110111,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m101000_0	),
Adb70100111000	(	adb70100111000,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m101000_0	),
Adb70100111001	(	adb70100111001,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m101000_0	),
Adb70100111010	(	adb70100111010,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m101000_0	),
Adb70100111011	(	adb70100111011,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m101000_0	),
Adb70100111100	(	adb70100111100,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m101000_0	),
Adb70100111101	(	adb70100111101,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m101000_0	),
Adb70100111110	(	adb70100111110,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m101000_0	),
Adb70100111111	(	adb70100111111,	n0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m101000_0	),
Adb70101000000	(	adb70101000000,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m101000_0	),
Adb70101000001	(	adb70101000001,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m101000_0	),
Adb70101000010	(	adb70101000010,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m101000_0	),
Adb70101000011	(	adb70101000011,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m101000_0	),
Adb70101000100	(	adb70101000100,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m101000_0	),
Adb70101000101	(	adb70101000101,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m101000_0	),
Adb70101000110	(	adb70101000110,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m101000_0	),
Adb70101000111	(	adb70101000111,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m101000_0	),
Adb70101001000	(	adb70101001000,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m101000_0	),
Adb70101001001	(	adb70101001001,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m101000_0	),
Adb70101001010	(	adb70101001010,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m101000_0	),
Adb70101001011	(	adb70101001011,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m101000_0	),
Adb70101001100	(	adb70101001100,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m101000_0	),
Adb70101001101	(	adb70101001101,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m101000_0	),
Adb70101001110	(	adb70101001110,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m101000_0	),
Adb70101001111	(	adb70101001111,	n0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m101000_0	),
Adb70101010000	(	adb70101010000,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m101000_0	),
Adb70101010001	(	adb70101010001,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m101000_0	),
Adb70101010010	(	adb70101010010,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m101000_0	),
Adb70101010011	(	adb70101010011,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m101000_0	),
Adb70101010100	(	adb70101010100,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m101000_0	),
Adb70101010101	(	adb70101010101,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m101000_0	),
Adb70101010110	(	adb70101010110,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m101000_0	),
Adb70101010111	(	adb70101010111,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m101000_0	),
Adb70101011000	(	adb70101011000,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m101000_0	),
Adb70101011001	(	adb70101011001,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m101000_0	),
Adb70101011010	(	adb70101011010,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m101000_0	),
Adb70101011011	(	adb70101011011,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m101000_0	),
Adb70101011100	(	adb70101011100,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m101000_0	),
Adb70101011101	(	adb70101011101,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m101000_0	),
Adb70101011110	(	adb70101011110,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m101000_0	),
Adb70101011111	(	adb70101011111,	n0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m101000_0	),
Adb70101100000	(	adb70101100000,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m101000_0	),
Adb70101100001	(	adb70101100001,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m101000_0	),
Adb70101100010	(	adb70101100010,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m101000_0	),
Adb70101100011	(	adb70101100011,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m101000_0	),
Adb70101100100	(	adb70101100100,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m101000_0	),
Adb70101100101	(	adb70101100101,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m101000_0	),
Adb70101100110	(	adb70101100110,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m101000_0	),
Adb70101100111	(	adb70101100111,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m101000_0	),
Adb70101101000	(	adb70101101000,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m101000_0	),
Adb70101101001	(	adb70101101001,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m101000_0	),
Adb70101101010	(	adb70101101010,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m101000_0	),
Adb70101101011	(	adb70101101011,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m101000_0	),
Adb70101101100	(	adb70101101100,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m101000_0	),
Adb70101101101	(	adb70101101101,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m101000_0	),
Adb70101101110	(	adb70101101110,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m101000_0	),
Adb70101101111	(	adb70101101111,	n0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m101000_0	),
Adb70101110000	(	adb70101110000,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m101000_0	),
Adb70101110001	(	adb70101110001,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m101000_0	),
Adb70101110010	(	adb70101110010,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m101000_0	),
Adb70101110011	(	adb70101110011,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m101000_0	),
Adb70101110100	(	adb70101110100,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m101000_0	),
Adb70101110101	(	adb70101110101,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m101000_0	),
Adb70101110110	(	adb70101110110,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m101000_0	),
Adb70101110111	(	adb70101110111,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m101000_0	),
Adb70101111000	(	adb70101111000,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m101000_0	),
Adb70101111001	(	adb70101111001,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m101000_0	),
Adb70101111010	(	adb70101111010,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m101000_0	),
Adb70101111011	(	adb70101111011,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m101000_0	),
Adb70101111100	(	adb70101111100,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m101000_0	),
Adb70101111101	(	adb70101111101,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m101000_0	),
Adb70101111110	(	adb70101111110,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m101000_0	),
Adb70101111111	(	adb70101111111,	n0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m101000_0	),
Adb70110000000	(	adb70110000000,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m100000_0	),
Adb70110000001	(	adb70110000001,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m100000_0	),
Adb70110000010	(	adb70110000010,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m100000_0	),
Adb70110000011	(	adb70110000011,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m100000_0	),
Adb70110000100	(	adb70110000100,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m100000_0	),
Adb70110000101	(	adb70110000101,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m100000_0	),
Adb70110000110	(	adb70110000110,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m100000_0	),
Adb70110000111	(	adb70110000111,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m100000_0	),
Adb70110001000	(	adb70110001000,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m100000_0	),
Adb70110001001	(	adb70110001001,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m100000_0	),
Adb70110001010	(	adb70110001010,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m100000_0	),
Adb70110001011	(	adb70110001011,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m100000_0	),
Adb70110001100	(	adb70110001100,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m100000_0	),
Adb70110001101	(	adb70110001101,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m100000_0	),
Adb70110001110	(	adb70110001110,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m100000_0	),
Adb70110001111	(	adb70110001111,	n0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m100000_0	),
Adb70110010000	(	adb70110010000,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m100000_0	),
Adb70110010001	(	adb70110010001,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m100000_0	),
Adb70110010010	(	adb70110010010,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m100000_0	),
Adb70110010011	(	adb70110010011,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m100000_0	),
Adb70110010100	(	adb70110010100,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m100000_0	),
Adb70110010101	(	adb70110010101,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m100000_0	),
Adb70110010110	(	adb70110010110,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m100000_0	),
Adb70110010111	(	adb70110010111,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m100000_0	),
Adb70110011000	(	adb70110011000,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m100000_0	),
Adb70110011001	(	adb70110011001,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m100000_0	),
Adb70110011010	(	adb70110011010,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m100000_0	),
Adb70110011011	(	adb70110011011,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m100000_0	),
Adb70110011100	(	adb70110011100,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m100000_0	),
Adb70110011101	(	adb70110011101,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m100000_0	),
Adb70110011110	(	adb70110011110,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m100000_0	),
Adb70110011111	(	adb70110011111,	n0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m100000_0	),
Adb70110100000	(	adb70110100000,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m100000_0	),
Adb70110100001	(	adb70110100001,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m100000_0	),
Adb70110100010	(	adb70110100010,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m100000_0	),
Adb70110100011	(	adb70110100011,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m100000_0	),
Adb70110100100	(	adb70110100100,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m100000_0	),
Adb70110100101	(	adb70110100101,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m100000_0	),
Adb70110100110	(	adb70110100110,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m100000_0	),
Adb70110100111	(	adb70110100111,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m100000_0	),
Adb70110101000	(	adb70110101000,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m100000_0	),
Adb70110101001	(	adb70110101001,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m100000_0	),
Adb70110101010	(	adb70110101010,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m100000_0	),
Adb70110101011	(	adb70110101011,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m100000_0	),
Adb70110101100	(	adb70110101100,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m100000_0	),
Adb70110101101	(	adb70110101101,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m100000_0	),
Adb70110101110	(	adb70110101110,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m100000_0	),
Adb70110101111	(	adb70110101111,	n0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m100000_0	),
Adb70110110000	(	adb70110110000,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m100000_0	),
Adb70110110001	(	adb70110110001,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m100000_0	),
Adb70110110010	(	adb70110110010,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m100000_0	),
Adb70110110011	(	adb70110110011,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m100000_0	),
Adb70110110100	(	adb70110110100,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m100000_0	),
Adb70110110101	(	adb70110110101,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m100000_0	),
Adb70110110110	(	adb70110110110,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m100000_0	),
Adb70110110111	(	adb70110110111,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m100000_0	),
Adb70110111000	(	adb70110111000,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m100000_0	),
Adb70110111001	(	adb70110111001,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m100000_0	),
Adb70110111010	(	adb70110111010,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m100000_0	),
Adb70110111011	(	adb70110111011,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m100000_0	),
Adb70110111100	(	adb70110111100,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m100000_0	),
Adb70110111101	(	adb70110111101,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m100000_0	),
Adb70110111110	(	adb70110111110,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m100000_0	),
Adb70110111111	(	adb70110111111,	n0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m100000_0	),
Adb70111000000	(	adb70111000000,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m100000_0	),
Adb70111000001	(	adb70111000001,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m100000_0	),
Adb70111000010	(	adb70111000010,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m100000_0	),
Adb70111000011	(	adb70111000011,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m100000_0	),
Adb70111000100	(	adb70111000100,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m100000_0	),
Adb70111000101	(	adb70111000101,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m100000_0	),
Adb70111000110	(	adb70111000110,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m100000_0	),
Adb70111000111	(	adb70111000111,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m100000_0	),
Adb70111001000	(	adb70111001000,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m100000_0	),
Adb70111001001	(	adb70111001001,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m100000_0	),
Adb70111001010	(	adb70111001010,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m100000_0	),
Adb70111001011	(	adb70111001011,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m100000_0	),
Adb70111001100	(	adb70111001100,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m100000_0	),
Adb70111001101	(	adb70111001101,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m100000_0	),
Adb70111001110	(	adb70111001110,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m100000_0	),
Adb70111001111	(	adb70111001111,	n0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m100000_0	),
Adb70111010000	(	adb70111010000,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m100000_0	),
Adb70111010001	(	adb70111010001,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m100000_0	),
Adb70111010010	(	adb70111010010,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m100000_0	),
Adb70111010011	(	adb70111010011,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m100000_0	),
Adb70111010100	(	adb70111010100,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m100000_0	),
Adb70111010101	(	adb70111010101,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m100000_0	),
Adb70111010110	(	adb70111010110,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m100000_0	),
Adb70111010111	(	adb70111010111,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m100000_0	),
Adb70111011000	(	adb70111011000,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m100000_0	),
Adb70111011001	(	adb70111011001,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m100000_0	),
Adb70111011010	(	adb70111011010,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m100000_0	),
Adb70111011011	(	adb70111011011,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m100000_0	),
Adb70111011100	(	adb70111011100,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m100000_0	),
Adb70111011101	(	adb70111011101,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m100000_0	),
Adb70111011110	(	adb70111011110,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m100000_0	),
Adb70111011111	(	adb70111011111,	n0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m100000_0	),
Adb70111100000	(	adb70111100000,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m100000_0	),
Adb70111100001	(	adb70111100001,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m100000_0	),
Adb70111100010	(	adb70111100010,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m100000_0	),
Adb70111100011	(	adb70111100011,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m100000_0	),
Adb70111100100	(	adb70111100100,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m100000_0	),
Adb70111100101	(	adb70111100101,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m100000_0	),
Adb70111100110	(	adb70111100110,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m100000_0	),
Adb70111100111	(	adb70111100111,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m100000_0	),
Adb70111101000	(	adb70111101000,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m100000_0	),
Adb70111101001	(	adb70111101001,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m100000_0	),
Adb70111101010	(	adb70111101010,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m100000_0	),
Adb70111101011	(	adb70111101011,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m100000_0	),
Adb70111101100	(	adb70111101100,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m100000_0	),
Adb70111101101	(	adb70111101101,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m100000_0	),
Adb70111101110	(	adb70111101110,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m100000_0	),
Adb70111101111	(	adb70111101111,	n0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m100000_0	),
Adb70111110000	(	adb70111110000,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m100000_0	),
Adb70111110001	(	adb70111110001,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m100000_0	),
Adb70111110010	(	adb70111110010,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m100000_0	),
Adb70111110011	(	adb70111110011,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m100000_0	),
Adb70111110100	(	adb70111110100,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m100000_0	),
Adb70111110101	(	adb70111110101,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m100000_0	),
Adb70111110110	(	adb70111110110,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m100000_0	),
Adb70111110111	(	adb70111110111,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m100000_0	),
Adb70111111000	(	adb70111111000,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m100000_0	),
Adb70111111001	(	adb70111111001,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m100000_0	),
Adb70111111010	(	adb70111111010,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m100000_0	),
Adb70111111011	(	adb70111111011,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m100000_0	),
Adb70111111100	(	adb70111111100,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m100000_0	),
Adb70111111101	(	adb70111111101,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m100000_0	),
Adb70111111110	(	adb70111111110,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m100000_0	),
Adb70111111111	(	adb70111111111,	n0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m100000_0	),
Adb71000000000	(	adb71000000000,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m011000_0	),
Adb71000000001	(	adb71000000001,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m011000_0	),
Adb71000000010	(	adb71000000010,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m011000_0	),
Adb71000000011	(	adb71000000011,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m011000_0	),
Adb71000000100	(	adb71000000100,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m011000_0	),
Adb71000000101	(	adb71000000101,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m011000_0	),
Adb71000000110	(	adb71000000110,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m011000_0	),
Adb71000000111	(	adb71000000111,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m011000_0	),
Adb71000001000	(	adb71000001000,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m011000_0	),
Adb71000001001	(	adb71000001001,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m011000_0	),
Adb71000001010	(	adb71000001010,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m011000_0	),
Adb71000001011	(	adb71000001011,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m011000_0	),
Adb71000001100	(	adb71000001100,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m011000_0	),
Adb71000001101	(	adb71000001101,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m011000_0	),
Adb71000001110	(	adb71000001110,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m011000_0	),
Adb71000001111	(	adb71000001111,	m0019,	n0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m011000_0	),
Adb71000010000	(	adb71000010000,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m011000_0	),
Adb71000010001	(	adb71000010001,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m011000_0	),
Adb71000010010	(	adb71000010010,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m011000_0	),
Adb71000010011	(	adb71000010011,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m011000_0	),
Adb71000010100	(	adb71000010100,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m011000_0	),
Adb71000010101	(	adb71000010101,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m011000_0	),
Adb71000010110	(	adb71000010110,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m011000_0	),
Adb71000010111	(	adb71000010111,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m011000_0	),
Adb71000011000	(	adb71000011000,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m011000_0	),
Adb71000011001	(	adb71000011001,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m011000_0	),
Adb71000011010	(	adb71000011010,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m011000_0	),
Adb71000011011	(	adb71000011011,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m011000_0	),
Adb71000011100	(	adb71000011100,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m011000_0	),
Adb71000011101	(	adb71000011101,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m011000_0	),
Adb71000011110	(	adb71000011110,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m011000_0	),
Adb71000011111	(	adb71000011111,	m0019,	n0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m011000_0	),
Adb71000100000	(	adb71000100000,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m011000_0	),
Adb71000100001	(	adb71000100001,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m011000_0	),
Adb71000100010	(	adb71000100010,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m011000_0	),
Adb71000100011	(	adb71000100011,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m011000_0	),
Adb71000100100	(	adb71000100100,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m011000_0	),
Adb71000100101	(	adb71000100101,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m011000_0	),
Adb71000100110	(	adb71000100110,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m011000_0	),
Adb71000100111	(	adb71000100111,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m011000_0	),
Adb71000101000	(	adb71000101000,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m011000_0	),
Adb71000101001	(	adb71000101001,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m011000_0	),
Adb71000101010	(	adb71000101010,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m011000_0	),
Adb71000101011	(	adb71000101011,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m011000_0	),
Adb71000101100	(	adb71000101100,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m011000_0	),
Adb71000101101	(	adb71000101101,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m011000_0	),
Adb71000101110	(	adb71000101110,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m011000_0	),
Adb71000101111	(	adb71000101111,	m0019,	n0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m011000_0	),
Adb71000110000	(	adb71000110000,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m011000_0	),
Adb71000110001	(	adb71000110001,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m011000_0	),
Adb71000110010	(	adb71000110010,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m011000_0	),
Adb71000110011	(	adb71000110011,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m011000_0	),
Adb71000110100	(	adb71000110100,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m011000_0	),
Adb71000110101	(	adb71000110101,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m011000_0	),
Adb71000110110	(	adb71000110110,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m011000_0	),
Adb71000110111	(	adb71000110111,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m011000_0	),
Adb71000111000	(	adb71000111000,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m011000_0	),
Adb71000111001	(	adb71000111001,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m011000_0	),
Adb71000111010	(	adb71000111010,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m011000_0	),
Adb71000111011	(	adb71000111011,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m011000_0	),
Adb71000111100	(	adb71000111100,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m011000_0	),
Adb71000111101	(	adb71000111101,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m011000_0	),
Adb71000111110	(	adb71000111110,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m011000_0	),
Adb71000111111	(	adb71000111111,	m0019,	n0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m011000_0	),
Adb71001000000	(	adb71001000000,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m011000_0	),
Adb71001000001	(	adb71001000001,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m011000_0	),
Adb71001000010	(	adb71001000010,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m011000_0	),
Adb71001000011	(	adb71001000011,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m011000_0	),
Adb71001000100	(	adb71001000100,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m011000_0	),
Adb71001000101	(	adb71001000101,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m011000_0	),
Adb71001000110	(	adb71001000110,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m011000_0	),
Adb71001000111	(	adb71001000111,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m011000_0	),
Adb71001001000	(	adb71001001000,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m011000_0	),
Adb71001001001	(	adb71001001001,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m011000_0	),
Adb71001001010	(	adb71001001010,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m011000_0	),
Adb71001001011	(	adb71001001011,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m011000_0	),
Adb71001001100	(	adb71001001100,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m011000_0	),
Adb71001001101	(	adb71001001101,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m011000_0	),
Adb71001001110	(	adb71001001110,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m011000_0	),
Adb71001001111	(	adb71001001111,	m0019,	n0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m011000_0	),
Adb71001010000	(	adb71001010000,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m011000_0	),
Adb71001010001	(	adb71001010001,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m011000_0	),
Adb71001010010	(	adb71001010010,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m011000_0	),
Adb71001010011	(	adb71001010011,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m011000_0	),
Adb71001010100	(	adb71001010100,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m011000_0	),
Adb71001010101	(	adb71001010101,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m011000_0	),
Adb71001010110	(	adb71001010110,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m011000_0	),
Adb71001010111	(	adb71001010111,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m011000_0	),
Adb71001011000	(	adb71001011000,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m011000_0	),
Adb71001011001	(	adb71001011001,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m011000_0	),
Adb71001011010	(	adb71001011010,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m011000_0	),
Adb71001011011	(	adb71001011011,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m011000_0	),
Adb71001011100	(	adb71001011100,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m011000_0	),
Adb71001011101	(	adb71001011101,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m011000_0	),
Adb71001011110	(	adb71001011110,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m011000_0	),
Adb71001011111	(	adb71001011111,	m0019,	n0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m011000_0	),
Adb71001100000	(	adb71001100000,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m011000_0	),
Adb71001100001	(	adb71001100001,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m011000_0	),
Adb71001100010	(	adb71001100010,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m011000_0	),
Adb71001100011	(	adb71001100011,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m011000_0	),
Adb71001100100	(	adb71001100100,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m011000_0	),
Adb71001100101	(	adb71001100101,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m011000_0	),
Adb71001100110	(	adb71001100110,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m011000_0	),
Adb71001100111	(	adb71001100111,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m011000_0	),
Adb71001101000	(	adb71001101000,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m011000_0	),
Adb71001101001	(	adb71001101001,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m011000_0	),
Adb71001101010	(	adb71001101010,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m011000_0	),
Adb71001101011	(	adb71001101011,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m011000_0	),
Adb71001101100	(	adb71001101100,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m011000_0	),
Adb71001101101	(	adb71001101101,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m011000_0	),
Adb71001101110	(	adb71001101110,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m011000_0	),
Adb71001101111	(	adb71001101111,	m0019,	n0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m011000_0	),
Adb71001110000	(	adb71001110000,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m011000_0	),
Adb71001110001	(	adb71001110001,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m011000_0	),
Adb71001110010	(	adb71001110010,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m011000_0	),
Adb71001110011	(	adb71001110011,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m011000_0	),
Adb71001110100	(	adb71001110100,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m011000_0	),
Adb71001110101	(	adb71001110101,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m011000_0	),
Adb71001110110	(	adb71001110110,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m011000_0	),
Adb71001110111	(	adb71001110111,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m011000_0	),
Adb71001111000	(	adb71001111000,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m011000_0	),
Adb71001111001	(	adb71001111001,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m011000_0	),
Adb71001111010	(	adb71001111010,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m011000_0	),
Adb71001111011	(	adb71001111011,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m011000_0	),
Adb71001111100	(	adb71001111100,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m011000_0	),
Adb71001111101	(	adb71001111101,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m011000_0	),
Adb71001111110	(	adb71001111110,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m011000_0	),
Adb71001111111	(	adb71001111111,	m0019,	n0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m011000_0	),
Adb71010000000	(	adb71010000000,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m010000_0	),
Adb71010000001	(	adb71010000001,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m010000_0	),
Adb71010000010	(	adb71010000010,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m010000_0	),
Adb71010000011	(	adb71010000011,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m010000_0	),
Adb71010000100	(	adb71010000100,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m010000_0	),
Adb71010000101	(	adb71010000101,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m010000_0	),
Adb71010000110	(	adb71010000110,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m010000_0	),
Adb71010000111	(	adb71010000111,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m010000_0	),
Adb71010001000	(	adb71010001000,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m010000_0	),
Adb71010001001	(	adb71010001001,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m010000_0	),
Adb71010001010	(	adb71010001010,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m010000_0	),
Adb71010001011	(	adb71010001011,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m010000_0	),
Adb71010001100	(	adb71010001100,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m010000_0	),
Adb71010001101	(	adb71010001101,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m010000_0	),
Adb71010001110	(	adb71010001110,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m010000_0	),
Adb71010001111	(	adb71010001111,	m0019,	n0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m010000_0	),
Adb71010010000	(	adb71010010000,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m010000_0	),
Adb71010010001	(	adb71010010001,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m010000_0	),
Adb71010010010	(	adb71010010010,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m010000_0	),
Adb71010010011	(	adb71010010011,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m010000_0	),
Adb71010010100	(	adb71010010100,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m010000_0	),
Adb71010010101	(	adb71010010101,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m010000_0	),
Adb71010010110	(	adb71010010110,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m010000_0	),
Adb71010010111	(	adb71010010111,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m010000_0	),
Adb71010011000	(	adb71010011000,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m010000_0	),
Adb71010011001	(	adb71010011001,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m010000_0	),
Adb71010011010	(	adb71010011010,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m010000_0	),
Adb71010011011	(	adb71010011011,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m010000_0	),
Adb71010011100	(	adb71010011100,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m010000_0	),
Adb71010011101	(	adb71010011101,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m010000_0	),
Adb71010011110	(	adb71010011110,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m010000_0	),
Adb71010011111	(	adb71010011111,	m0019,	n0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m010000_0	),
Adb71010100000	(	adb71010100000,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m010000_0	),
Adb71010100001	(	adb71010100001,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m010000_0	),
Adb71010100010	(	adb71010100010,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m010000_0	),
Adb71010100011	(	adb71010100011,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m010000_0	),
Adb71010100100	(	adb71010100100,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m010000_0	),
Adb71010100101	(	adb71010100101,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m010000_0	),
Adb71010100110	(	adb71010100110,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m010000_0	),
Adb71010100111	(	adb71010100111,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m010000_0	),
Adb71010101000	(	adb71010101000,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m010000_0	),
Adb71010101001	(	adb71010101001,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m010000_0	),
Adb71010101010	(	adb71010101010,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m010000_0	),
Adb71010101011	(	adb71010101011,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m010000_0	),
Adb71010101100	(	adb71010101100,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m010000_0	),
Adb71010101101	(	adb71010101101,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m010000_0	),
Adb71010101110	(	adb71010101110,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m010000_0	),
Adb71010101111	(	adb71010101111,	m0019,	n0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m010000_0	),
Adb71010110000	(	adb71010110000,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m010000_0	),
Adb71010110001	(	adb71010110001,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m010000_0	),
Adb71010110010	(	adb71010110010,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m010000_0	),
Adb71010110011	(	adb71010110011,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m010000_0	),
Adb71010110100	(	adb71010110100,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m010000_0	),
Adb71010110101	(	adb71010110101,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m010000_0	),
Adb71010110110	(	adb71010110110,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m010000_0	),
Adb71010110111	(	adb71010110111,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m010000_0	),
Adb71010111000	(	adb71010111000,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m010000_0	),
Adb71010111001	(	adb71010111001,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m010000_0	),
Adb71010111010	(	adb71010111010,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m010000_0	),
Adb71010111011	(	adb71010111011,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m010000_0	),
Adb71010111100	(	adb71010111100,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m010000_0	),
Adb71010111101	(	adb71010111101,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m010000_0	),
Adb71010111110	(	adb71010111110,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m010000_0	),
Adb71010111111	(	adb71010111111,	m0019,	n0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m010000_0	),
Adb71011000000	(	adb71011000000,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m010000_0	),
Adb71011000001	(	adb71011000001,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m010000_0	),
Adb71011000010	(	adb71011000010,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m010000_0	),
Adb71011000011	(	adb71011000011,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m010000_0	),
Adb71011000100	(	adb71011000100,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m010000_0	),
Adb71011000101	(	adb71011000101,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m010000_0	),
Adb71011000110	(	adb71011000110,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m010000_0	),
Adb71011000111	(	adb71011000111,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m010000_0	),
Adb71011001000	(	adb71011001000,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m010000_0	),
Adb71011001001	(	adb71011001001,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m010000_0	),
Adb71011001010	(	adb71011001010,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m010000_0	),
Adb71011001011	(	adb71011001011,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m010000_0	),
Adb71011001100	(	adb71011001100,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m010000_0	),
Adb71011001101	(	adb71011001101,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m010000_0	),
Adb71011001110	(	adb71011001110,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m010000_0	),
Adb71011001111	(	adb71011001111,	m0019,	n0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m010000_0	),
Adb71011010000	(	adb71011010000,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m010000_0	),
Adb71011010001	(	adb71011010001,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m010000_0	),
Adb71011010010	(	adb71011010010,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m010000_0	),
Adb71011010011	(	adb71011010011,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m010000_0	),
Adb71011010100	(	adb71011010100,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m010000_0	),
Adb71011010101	(	adb71011010101,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m010000_0	),
Adb71011010110	(	adb71011010110,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m010000_0	),
Adb71011010111	(	adb71011010111,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m010000_0	),
Adb71011011000	(	adb71011011000,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m010000_0	),
Adb71011011001	(	adb71011011001,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m010000_0	),
Adb71011011010	(	adb71011011010,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m010000_0	),
Adb71011011011	(	adb71011011011,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m010000_0	),
Adb71011011100	(	adb71011011100,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m010000_0	),
Adb71011011101	(	adb71011011101,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m010000_0	),
Adb71011011110	(	adb71011011110,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m010000_0	),
Adb71011011111	(	adb71011011111,	m0019,	n0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m010000_0	),
Adb71011100000	(	adb71011100000,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m010000_0	),
Adb71011100001	(	adb71011100001,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m010000_0	),
Adb71011100010	(	adb71011100010,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m010000_0	),
Adb71011100011	(	adb71011100011,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m010000_0	),
Adb71011100100	(	adb71011100100,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m010000_0	),
Adb71011100101	(	adb71011100101,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m010000_0	),
Adb71011100110	(	adb71011100110,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m010000_0	),
Adb71011100111	(	adb71011100111,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m010000_0	),
Adb71011101000	(	adb71011101000,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m010000_0	),
Adb71011101001	(	adb71011101001,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m010000_0	),
Adb71011101010	(	adb71011101010,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m010000_0	),
Adb71011101011	(	adb71011101011,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m010000_0	),
Adb71011101100	(	adb71011101100,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m010000_0	),
Adb71011101101	(	adb71011101101,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m010000_0	),
Adb71011101110	(	adb71011101110,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m010000_0	),
Adb71011101111	(	adb71011101111,	m0019,	n0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m010000_0	),
Adb71011110000	(	adb71011110000,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m010000_0	),
Adb71011110001	(	adb71011110001,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m010000_0	),
Adb71011110010	(	adb71011110010,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m010000_0	),
Adb71011110011	(	adb71011110011,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m010000_0	),
Adb71011110100	(	adb71011110100,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m010000_0	),
Adb71011110101	(	adb71011110101,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m010000_0	),
Adb71011110110	(	adb71011110110,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m010000_0	),
Adb71011110111	(	adb71011110111,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m010000_0	),
Adb71011111000	(	adb71011111000,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m010000_0	),
Adb71011111001	(	adb71011111001,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m010000_0	),
Adb71011111010	(	adb71011111010,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m010000_0	),
Adb71011111011	(	adb71011111011,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m010000_0	),
Adb71011111100	(	adb71011111100,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m010000_0	),
Adb71011111101	(	adb71011111101,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m010000_0	),
Adb71011111110	(	adb71011111110,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m010000_0	),
Adb71011111111	(	adb71011111111,	m0019,	n0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m010000_0	),
Adb71100000000	(	adb71100000000,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m001000_0	),
Adb71100000001	(	adb71100000001,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m001000_0	),
Adb71100000010	(	adb71100000010,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m001000_0	),
Adb71100000011	(	adb71100000011,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m001000_0	),
Adb71100000100	(	adb71100000100,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m001000_0	),
Adb71100000101	(	adb71100000101,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m001000_0	),
Adb71100000110	(	adb71100000110,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m001000_0	),
Adb71100000111	(	adb71100000111,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m001000_0	),
Adb71100001000	(	adb71100001000,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m001000_0	),
Adb71100001001	(	adb71100001001,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m001000_0	),
Adb71100001010	(	adb71100001010,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m001000_0	),
Adb71100001011	(	adb71100001011,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m001000_0	),
Adb71100001100	(	adb71100001100,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m001000_0	),
Adb71100001101	(	adb71100001101,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m001000_0	),
Adb71100001110	(	adb71100001110,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m001000_0	),
Adb71100001111	(	adb71100001111,	m0019,	m0018,	n0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m001000_0	),
Adb71100010000	(	adb71100010000,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m001000_0	),
Adb71100010001	(	adb71100010001,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m001000_0	),
Adb71100010010	(	adb71100010010,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m001000_0	),
Adb71100010011	(	adb71100010011,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m001000_0	),
Adb71100010100	(	adb71100010100,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m001000_0	),
Adb71100010101	(	adb71100010101,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m001000_0	),
Adb71100010110	(	adb71100010110,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m001000_0	),
Adb71100010111	(	adb71100010111,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m001000_0	),
Adb71100011000	(	adb71100011000,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m001000_0	),
Adb71100011001	(	adb71100011001,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m001000_0	),
Adb71100011010	(	adb71100011010,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m001000_0	),
Adb71100011011	(	adb71100011011,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m001000_0	),
Adb71100011100	(	adb71100011100,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m001000_0	),
Adb71100011101	(	adb71100011101,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m001000_0	),
Adb71100011110	(	adb71100011110,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m001000_0	),
Adb71100011111	(	adb71100011111,	m0019,	m0018,	n0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m001000_0	),
Adb71100100000	(	adb71100100000,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m001000_0	),
Adb71100100001	(	adb71100100001,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m001000_0	),
Adb71100100010	(	adb71100100010,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m001000_0	),
Adb71100100011	(	adb71100100011,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m001000_0	),
Adb71100100100	(	adb71100100100,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m001000_0	),
Adb71100100101	(	adb71100100101,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m001000_0	),
Adb71100100110	(	adb71100100110,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m001000_0	),
Adb71100100111	(	adb71100100111,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m001000_0	),
Adb71100101000	(	adb71100101000,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m001000_0	),
Adb71100101001	(	adb71100101001,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m001000_0	),
Adb71100101010	(	adb71100101010,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m001000_0	),
Adb71100101011	(	adb71100101011,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m001000_0	),
Adb71100101100	(	adb71100101100,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m001000_0	),
Adb71100101101	(	adb71100101101,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m001000_0	),
Adb71100101110	(	adb71100101110,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m001000_0	),
Adb71100101111	(	adb71100101111,	m0019,	m0018,	n0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m001000_0	),
Adb71100110000	(	adb71100110000,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m001000_0	),
Adb71100110001	(	adb71100110001,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m001000_0	),
Adb71100110010	(	adb71100110010,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m001000_0	),
Adb71100110011	(	adb71100110011,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m001000_0	),
Adb71100110100	(	adb71100110100,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m001000_0	),
Adb71100110101	(	adb71100110101,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m001000_0	),
Adb71100110110	(	adb71100110110,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m001000_0	),
Adb71100110111	(	adb71100110111,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m001000_0	),
Adb71100111000	(	adb71100111000,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m001000_0	),
Adb71100111001	(	adb71100111001,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m001000_0	),
Adb71100111010	(	adb71100111010,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m001000_0	),
Adb71100111011	(	adb71100111011,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m001000_0	),
Adb71100111100	(	adb71100111100,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m001000_0	),
Adb71100111101	(	adb71100111101,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m001000_0	),
Adb71100111110	(	adb71100111110,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m001000_0	),
Adb71100111111	(	adb71100111111,	m0019,	m0018,	n0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m001000_0	),
Adb71101000000	(	adb71101000000,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m001000_0	),
Adb71101000001	(	adb71101000001,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m001000_0	),
Adb71101000010	(	adb71101000010,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m001000_0	),
Adb71101000011	(	adb71101000011,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m001000_0	),
Adb71101000100	(	adb71101000100,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m001000_0	),
Adb71101000101	(	adb71101000101,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m001000_0	),
Adb71101000110	(	adb71101000110,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m001000_0	),
Adb71101000111	(	adb71101000111,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m001000_0	),
Adb71101001000	(	adb71101001000,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m001000_0	),
Adb71101001001	(	adb71101001001,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m001000_0	),
Adb71101001010	(	adb71101001010,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m001000_0	),
Adb71101001011	(	adb71101001011,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m001000_0	),
Adb71101001100	(	adb71101001100,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m001000_0	),
Adb71101001101	(	adb71101001101,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m001000_0	),
Adb71101001110	(	adb71101001110,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m001000_0	),
Adb71101001111	(	adb71101001111,	m0019,	m0018,	n0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m001000_0	),
Adb71101010000	(	adb71101010000,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m001000_0	),
Adb71101010001	(	adb71101010001,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m001000_0	),
Adb71101010010	(	adb71101010010,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m001000_0	),
Adb71101010011	(	adb71101010011,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m001000_0	),
Adb71101010100	(	adb71101010100,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m001000_0	),
Adb71101010101	(	adb71101010101,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m001000_0	),
Adb71101010110	(	adb71101010110,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m001000_0	),
Adb71101010111	(	adb71101010111,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m001000_0	),
Adb71101011000	(	adb71101011000,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m001000_0	),
Adb71101011001	(	adb71101011001,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m001000_0	),
Adb71101011010	(	adb71101011010,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m001000_0	),
Adb71101011011	(	adb71101011011,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m001000_0	),
Adb71101011100	(	adb71101011100,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m001000_0	),
Adb71101011101	(	adb71101011101,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m001000_0	),
Adb71101011110	(	adb71101011110,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m001000_0	),
Adb71101011111	(	adb71101011111,	m0019,	m0018,	n0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m001000_0	),
Adb71101100000	(	adb71101100000,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m001000_0	),
Adb71101100001	(	adb71101100001,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m001000_0	),
Adb71101100010	(	adb71101100010,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m001000_0	),
Adb71101100011	(	adb71101100011,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m001000_0	),
Adb71101100100	(	adb71101100100,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m001000_0	),
Adb71101100101	(	adb71101100101,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m001000_0	),
Adb71101100110	(	adb71101100110,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m001000_0	),
Adb71101100111	(	adb71101100111,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m001000_0	),
Adb71101101000	(	adb71101101000,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m001000_0	),
Adb71101101001	(	adb71101101001,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m001000_0	),
Adb71101101010	(	adb71101101010,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m001000_0	),
Adb71101101011	(	adb71101101011,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m001000_0	),
Adb71101101100	(	adb71101101100,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m001000_0	),
Adb71101101101	(	adb71101101101,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m001000_0	),
Adb71101101110	(	adb71101101110,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m001000_0	),
Adb71101101111	(	adb71101101111,	m0019,	m0018,	n0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m001000_0	),
Adb71101110000	(	adb71101110000,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m001000_0	),
Adb71101110001	(	adb71101110001,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m001000_0	),
Adb71101110010	(	adb71101110010,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m001000_0	),
Adb71101110011	(	adb71101110011,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m001000_0	),
Adb71101110100	(	adb71101110100,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m001000_0	),
Adb71101110101	(	adb71101110101,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m001000_0	),
Adb71101110110	(	adb71101110110,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m001000_0	),
Adb71101110111	(	adb71101110111,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m001000_0	),
Adb71101111000	(	adb71101111000,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m001000_0	),
Adb71101111001	(	adb71101111001,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m001000_0	),
Adb71101111010	(	adb71101111010,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m001000_0	),
Adb71101111011	(	adb71101111011,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m001000_0	),
Adb71101111100	(	adb71101111100,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m001000_0	),
Adb71101111101	(	adb71101111101,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m001000_0	),
Adb71101111110	(	adb71101111110,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m001000_0	),
Adb71101111111	(	adb71101111111,	m0019,	m0018,	n0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m001000_0	),
Adb71110000000	(	adb71110000000,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0000000_0,	m000000_0	),
Adb71110000001	(	adb71110000001,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0000001_0,	m000000_0	),
Adb71110000010	(	adb71110000010,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0000010_0,	m000000_0	),
Adb71110000011	(	adb71110000011,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0000011_0,	m000000_0	),
Adb71110000100	(	adb71110000100,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0000100_0,	m000000_0	),
Adb71110000101	(	adb71110000101,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0000101_0,	m000000_0	),
Adb71110000110	(	adb71110000110,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0000110_0,	m000000_0	),
Adb71110000111	(	adb71110000111,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0000111_0,	m000000_0	),
Adb71110001000	(	adb71110001000,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0001000_0,	m000000_0	),
Adb71110001001	(	adb71110001001,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0001001_0,	m000000_0	),
Adb71110001010	(	adb71110001010,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0001010_0,	m000000_0	),
Adb71110001011	(	adb71110001011,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0001011_0,	m000000_0	),
Adb71110001100	(	adb71110001100,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0001100_0,	m000000_0	),
Adb71110001101	(	adb71110001101,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0001101_0,	m000000_0	),
Adb71110001110	(	adb71110001110,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0001110_0,	m000000_0	),
Adb71110001111	(	adb71110001111,	m0019,	m0018,	m0017,	n0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0001111_0,	m000000_0	),
Adb71110010000	(	adb71110010000,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0010000_0,	m000000_0	),
Adb71110010001	(	adb71110010001,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0010001_0,	m000000_0	),
Adb71110010010	(	adb71110010010,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0010010_0,	m000000_0	),
Adb71110010011	(	adb71110010011,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0010011_0,	m000000_0	),
Adb71110010100	(	adb71110010100,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0010100_0,	m000000_0	),
Adb71110010101	(	adb71110010101,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0010101_0,	m000000_0	),
Adb71110010110	(	adb71110010110,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0010110_0,	m000000_0	),
Adb71110010111	(	adb71110010111,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0010111_0,	m000000_0	),
Adb71110011000	(	adb71110011000,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0011000_0,	m000000_0	),
Adb71110011001	(	adb71110011001,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0011001_0,	m000000_0	),
Adb71110011010	(	adb71110011010,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0011010_0,	m000000_0	),
Adb71110011011	(	adb71110011011,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0011011_0,	m000000_0	),
Adb71110011100	(	adb71110011100,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0011100_0,	m000000_0	),
Adb71110011101	(	adb71110011101,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0011101_0,	m000000_0	),
Adb71110011110	(	adb71110011110,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0011110_0,	m000000_0	),
Adb71110011111	(	adb71110011111,	m0019,	m0018,	m0017,	n0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0011111_0,	m000000_0	),
Adb71110100000	(	adb71110100000,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0100000_0,	m000000_0	),
Adb71110100001	(	adb71110100001,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0100001_0,	m000000_0	),
Adb71110100010	(	adb71110100010,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0100010_0,	m000000_0	),
Adb71110100011	(	adb71110100011,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0100011_0,	m000000_0	),
Adb71110100100	(	adb71110100100,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0100100_0,	m000000_0	),
Adb71110100101	(	adb71110100101,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0100101_0,	m000000_0	),
Adb71110100110	(	adb71110100110,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0100110_0,	m000000_0	),
Adb71110100111	(	adb71110100111,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0100111_0,	m000000_0	),
Adb71110101000	(	adb71110101000,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0101000_0,	m000000_0	),
Adb71110101001	(	adb71110101001,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0101001_0,	m000000_0	),
Adb71110101010	(	adb71110101010,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0101010_0,	m000000_0	),
Adb71110101011	(	adb71110101011,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0101011_0,	m000000_0	),
Adb71110101100	(	adb71110101100,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0101100_0,	m000000_0	),
Adb71110101101	(	adb71110101101,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0101101_0,	m000000_0	),
Adb71110101110	(	adb71110101110,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0101110_0,	m000000_0	),
Adb71110101111	(	adb71110101111,	m0019,	m0018,	m0017,	n0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0101111_0,	m000000_0	),
Adb71110110000	(	adb71110110000,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m0110000_0,	m000000_0	),
Adb71110110001	(	adb71110110001,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m0110001_0,	m000000_0	),
Adb71110110010	(	adb71110110010,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m0110010_0,	m000000_0	),
Adb71110110011	(	adb71110110011,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m0110011_0,	m000000_0	),
Adb71110110100	(	adb71110110100,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m0110100_0,	m000000_0	),
Adb71110110101	(	adb71110110101,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m0110101_0,	m000000_0	),
Adb71110110110	(	adb71110110110,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m0110110_0,	m000000_0	),
Adb71110110111	(	adb71110110111,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m0110111_0,	m000000_0	),
Adb71110111000	(	adb71110111000,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m0111000_0,	m000000_0	),
Adb71110111001	(	adb71110111001,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m0111001_0,	m000000_0	),
Adb71110111010	(	adb71110111010,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m0111010_0,	m000000_0	),
Adb71110111011	(	adb71110111011,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m0111011_0,	m000000_0	),
Adb71110111100	(	adb71110111100,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m0111100_0,	m000000_0	),
Adb71110111101	(	adb71110111101,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m0111101_0,	m000000_0	),
Adb71110111110	(	adb71110111110,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m0111110_0,	m000000_0	),
Adb71110111111	(	adb71110111111,	m0019,	m0018,	m0017,	n0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m0111111_0,	m000000_0	),
Adb71111000000	(	adb71111000000,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1000000_0,	m000000_0	),
Adb71111000001	(	adb71111000001,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1000001_0,	m000000_0	),
Adb71111000010	(	adb71111000010,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1000010_0,	m000000_0	),
Adb71111000011	(	adb71111000011,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1000011_0,	m000000_0	),
Adb71111000100	(	adb71111000100,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1000100_0,	m000000_0	),
Adb71111000101	(	adb71111000101,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1000101_0,	m000000_0	),
Adb71111000110	(	adb71111000110,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1000110_0,	m000000_0	),
Adb71111000111	(	adb71111000111,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1000111_0,	m000000_0	),
Adb71111001000	(	adb71111001000,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1001000_0,	m000000_0	),
Adb71111001001	(	adb71111001001,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1001001_0,	m000000_0	),
Adb71111001010	(	adb71111001010,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1001010_0,	m000000_0	),
Adb71111001011	(	adb71111001011,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1001011_0,	m000000_0	),
Adb71111001100	(	adb71111001100,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1001100_0,	m000000_0	),
Adb71111001101	(	adb71111001101,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1001101_0,	m000000_0	),
Adb71111001110	(	adb71111001110,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1001110_0,	m000000_0	),
Adb71111001111	(	adb71111001111,	m0019,	m0018,	m0017,	m0016,	n0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1001111_0,	m000000_0	),
Adb71111010000	(	adb71111010000,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1010000_0,	m000000_0	),
Adb71111010001	(	adb71111010001,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1010001_0,	m000000_0	),
Adb71111010010	(	adb71111010010,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1010010_0,	m000000_0	),
Adb71111010011	(	adb71111010011,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1010011_0,	m000000_0	),
Adb71111010100	(	adb71111010100,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1010100_0,	m000000_0	),
Adb71111010101	(	adb71111010101,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1010101_0,	m000000_0	),
Adb71111010110	(	adb71111010110,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1010110_0,	m000000_0	),
Adb71111010111	(	adb71111010111,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1010111_0,	m000000_0	),
Adb71111011000	(	adb71111011000,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1011000_0,	m000000_0	),
Adb71111011001	(	adb71111011001,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1011001_0,	m000000_0	),
Adb71111011010	(	adb71111011010,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1011010_0,	m000000_0	),
Adb71111011011	(	adb71111011011,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1011011_0,	m000000_0	),
Adb71111011100	(	adb71111011100,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1011100_0,	m000000_0	),
Adb71111011101	(	adb71111011101,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1011101_0,	m000000_0	),
Adb71111011110	(	adb71111011110,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1011110_0,	m000000_0	),
Adb71111011111	(	adb71111011111,	m0019,	m0018,	m0017,	m0016,	n0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1011111_0,	m000000_0	),
Adb71111100000	(	adb71111100000,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1100000_0,	m000000_0	),
Adb71111100001	(	adb71111100001,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1100001_0,	m000000_0	),
Adb71111100010	(	adb71111100010,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1100010_0,	m000000_0	),
Adb71111100011	(	adb71111100011,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1100011_0,	m000000_0	),
Adb71111100100	(	adb71111100100,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1100100_0,	m000000_0	),
Adb71111100101	(	adb71111100101,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1100101_0,	m000000_0	),
Adb71111100110	(	adb71111100110,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1100110_0,	m000000_0	),
Adb71111100111	(	adb71111100111,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1100111_0,	m000000_0	),
Adb71111101000	(	adb71111101000,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1101000_0,	m000000_0	),
Adb71111101001	(	adb71111101001,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1101001_0,	m000000_0	),
Adb71111101010	(	adb71111101010,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1101010_0,	m000000_0	),
Adb71111101011	(	adb71111101011,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1101011_0,	m000000_0	),
Adb71111101100	(	adb71111101100,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1101100_0,	m000000_0	),
Adb71111101101	(	adb71111101101,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1101101_0,	m000000_0	),
Adb71111101110	(	adb71111101110,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1101110_0,	m000000_0	),
Adb71111101111	(	adb71111101111,	m0019,	m0018,	m0017,	m0016,	m0015,	n0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1101111_0,	m000000_0	),
Adb71111110000	(	adb71111110000,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	n0009,	m1110000_0,	m000000_0	),
Adb71111110001	(	adb71111110001,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	n0010,	m0009,	m1110001_0,	m000000_0	),
Adb71111110010	(	adb71111110010,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	n0009,	m1110010_0,	m000000_0	),
Adb71111110011	(	adb71111110011,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	n0012,	m0011,	m0010,	m0009,	m1110011_0,	m000000_0	),
Adb71111110100	(	adb71111110100,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	n0009,	m1110100_0,	m000000_0	),
Adb71111110101	(	adb71111110101,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	n0010,	m0009,	m1110101_0,	m000000_0	),
Adb71111110110	(	adb71111110110,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	n0009,	m1110110_0,	m000000_0	),
Adb71111110111	(	adb71111110111,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	n0013,	m0012,	m0011,	m0010,	m0009,	m1110111_0,	m000000_0	),
Adb71111111000	(	adb71111111000,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	n0009,	m1111000_0,	m000000_0	),
Adb71111111001	(	adb71111111001,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	n0010,	m0009,	m1111001_0,	m000000_0	),
Adb71111111010	(	adb71111111010,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	n0009,	m1111010_0,	m000000_0	),
Adb71111111011	(	adb71111111011,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	n0012,	m0011,	m0010,	m0009,	m1111011_0,	m000000_0	),
Adb71111111100	(	adb71111111100,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	n0009,	m1111100_0,	m000000_0	),
Adb71111111101	(	adb71111111101,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	n0010,	m0009,	m1111101_0,	m000000_0	),
Adb71111111110	(	adb71111111110,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	n0009,	m1111110_0,	m000000_0	),
Adb71111111111	(	adb71111111111,	m0019,	m0018,	m0017,	m0016,	m0015,	m0014,	m0013,	m0012,	m0011,	m0010,	m0009,	m1111111_0,	m000000_0	),
       Adbtopline0(adbtopline0,n0019,n0018,n0017,m0011),
       Adbtopline1(adbtopline1,m0019,m0018,m0017,m0011),
       Adbp102(adbp102,m0019,m0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m102_0),
       Adbp103(adbp103,m0019,m0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m103_0),
       Adbp104(adbp104,m0019,m0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m104_0),
       Adbp105(adbp105,m0019,m0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m105_0),
       Adbp106(adbp106,m0019,m0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m106_0),
       Adbp107(adbp107,m0019,m0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m107_0),
       Adbp108(adbp108,m0019,m0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m108_0),
       Adbp109(adbp109,m0019,m0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m109_0),
       Adbp110(adbp110,m0019,m0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m110_0),
       Adbp111(adbp111,m0019,m0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m111_0),
       Adbp112(adbp112,m0019,m0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m112_0),
       Adbp113(adbp113,m0019,m0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m113_0),
       Adbp114(adbp114,m0019,m0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m114_0),
       Adbp115(adbp115,m0019,m0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m115_0),
       Adbp116(adbp116,m0019,n0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m116_0),
       Adbp117(adbp117,m0019,n0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m117_0),
       Adbp118(adbp118,m0019,n0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m118_0),
       Adbp119(adbp119,m0019,n0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m119_0),
       Adbp120(adbp120,m0019,n0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m120_0),
       Adbp121(adbp121,m0019,n0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m121_0),
       Adbp122(adbp122,m0019,n0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m122_0),
       Adbp123(adbp123,m0019,n0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m123_0),
       Adbp124(adbp124,m0019,n0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m124_0),
       Adbp125(adbp125,m0019,n0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m125_0),
       Adbp126(adbp126,m0019,n0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m126_0),
       Adbp127(adbp127,m0019,n0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m127_0),
       Adbp128(adbp128,m0019,n0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m128_0),
       Adbp129(adbp129,m0019,n0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m129_0),
       Adbp130(adbp130,m0019,n0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m130_0),
       Adbp131(adbp131,m0019,n0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m131_0),
       Adbp132(adbp132,n0019,m0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m132_0),
       Adbp133(adbp133,n0019,m0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m133_0),
       Adbp134(adbp134,n0019,m0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m134_0),
       Adbp135(adbp135,n0019,m0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m135_0),
       Adbp136(adbp136,n0019,m0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m136_0),
       Adbp137(adbp137,n0019,m0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m137_0),
       Adbp138(adbp138,n0019,m0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m138_0),
       Adbp139(adbp139,n0019,m0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m139_0),
       Adbp140(adbp140,n0019,m0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m140_0),
       Adbp141(adbp141,n0019,m0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m141_0),
       Adbp142(adbp142,n0019,m0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m142_0),
       Adbp143(adbp143,n0019,m0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m143_0),
       Adbp144(adbp144,n0019,m0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m144_0),
       Adbp145(adbp145,n0019,m0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m145_0),
       Adbp146(adbp146,n0019,m0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m146_0),
       Adbp147(adbp147,n0019,m0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m147_0),
       Adbp148(adbp148,n0019,n0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m148_0),
       Adbp149(adbp149,n0019,n0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m149_0),
       Adbp150(adbp150,n0019,n0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m150_0),
       Adbp151(adbp151,n0019,n0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m151_0),
       Adbp152(adbp152,n0019,n0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m152_0),
       Adbp153(adbp153,n0019,n0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m153_0),
       Adbp154(adbp154,n0019,n0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m154_0),
       Adbp155(adbp155,n0019,n0018,m0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m155_0),
       Adbp156(adbp156,n0019,n0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m156_0),
       Adbp157(adbp157,n0019,n0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m157_0),
       Adbp158(adbp158,n0019,n0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m158_0),
       Adbp159(adbp159,n0019,n0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m159_0),
       Adbp160(adbp160,n0019,n0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m160_0),
       Adbp161(adbp161,n0019,n0018,n0017,n0016,n0015,n0014,n0013,m0012,m0011,n0010,m161_0),
       Adbp202(adbp202,m0019,m0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m202_0),
       Adbp203(adbp203,m0019,m0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m203_0),
       Adbp204(adbp204,m0019,m0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m204_0),
       Adbp205(adbp205,m0019,m0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m205_0),
       Adbp206(adbp206,m0019,m0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m206_0),
       Adbp207(adbp207,m0019,m0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m207_0),
       Adbp208(adbp208,m0019,m0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m208_0),
       Adbp209(adbp209,m0019,m0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m209_0),
       Adbp210(adbp210,m0019,m0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m210_0),
       Adbp211(adbp211,m0019,m0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m211_0),
       Adbp212(adbp212,m0019,m0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m212_0),
       Adbp213(adbp213,m0019,m0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m213_0),
       Adbp214(adbp214,m0019,m0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m214_0),
       Adbp215(adbp215,m0019,m0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m215_0),
       Adbp216(adbp216,m0019,n0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m216_0),
       Adbp217(adbp217,m0019,n0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m217_0),
       Adbp218(adbp218,m0019,n0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m218_0),
       Adbp219(adbp219,m0019,n0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m219_0),
       Adbp220(adbp220,m0019,n0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m220_0),
       Adbp221(adbp221,m0019,n0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m221_0),
       Adbp222(adbp222,m0019,n0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m222_0),
       Adbp223(adbp223,m0019,n0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m223_0),
       Adbp224(adbp224,m0019,n0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m224_0),
       Adbp225(adbp225,m0019,n0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m225_0),
       Adbp226(adbp226,m0019,n0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m226_0),
       Adbp227(adbp227,m0019,n0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m227_0),
       Adbp228(adbp228,m0019,n0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m228_0),
       Adbp229(adbp229,m0019,n0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m229_0),
       Adbp230(adbp230,m0019,n0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m230_0),
       Adbp231(adbp231,m0019,n0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m231_0),
       Adbp232(adbp232,n0019,m0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m232_0),
       Adbp233(adbp233,n0019,m0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m233_0),
       Adbp234(adbp234,n0019,m0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m234_0),
       Adbp235(adbp235,n0019,m0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m235_0),
       Adbp236(adbp236,n0019,m0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m236_0),
       Adbp237(adbp237,n0019,m0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m237_0),
       Adbp238(adbp238,n0019,m0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m238_0),
       Adbp239(adbp239,n0019,m0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m239_0),
       Adbp240(adbp240,n0019,m0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m240_0),
       Adbp241(adbp241,n0019,m0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m241_0),
       Adbp242(adbp242,n0019,m0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m242_0),
       Adbp243(adbp243,n0019,m0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m243_0),
       Adbp244(adbp244,n0019,m0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m244_0),
       Adbp245(adbp245,n0019,m0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m245_0),
       Adbp246(adbp246,n0019,m0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m246_0),
       Adbp247(adbp247,n0019,m0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m247_0),
       Adbp248(adbp248,n0019,n0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m248_0),
       Adbp249(adbp249,n0019,n0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m249_0),
       Adbp250(adbp250,n0019,n0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m250_0),
       Adbp251(adbp251,n0019,n0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m251_0),
       Adbp252(adbp252,n0019,n0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m252_0),
       Adbp253(adbp253,n0019,n0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m253_0),
       Adbp254(adbp254,n0019,n0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m254_0),
       Adbp255(adbp255,n0019,n0018,m0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m255_0),
       Adbp256(adbp256,n0019,n0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m256_0),
       Adbp257(adbp257,n0019,n0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m257_0),
       Adbp258(adbp258,n0019,n0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m258_0),
       Adbp259(adbp259,n0019,n0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m259_0),
       Adbp260(adbp260,n0019,n0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m260_0),
       Adbp261(adbp261,n0019,n0018,n0017,m0016,m0015,m0014,m0013,n0012,m0011,m0010,m261_0);

initial begin
m0000000_0=0;
q0000000_0=0;
m0000000_1=0;
q0000000_1=0;
m0000001_0=0;
q0000001_0=0;
m0000001_1=0;
q0000001_1=0;
m0000010_0=0;
q0000010_0=0;
m0000010_1=0;
q0000010_1=0;
m0000011_0=0;
q0000011_0=0;
m0000011_1=0;
q0000011_1=0;
m0000100_0=0;
q0000100_0=0;
m0000100_1=0;
q0000100_1=0;
m0000101_0=0;
q0000101_0=0;
m0000101_1=0;
q0000101_1=0;
m0000110_0=0;
q0000110_0=0;
m0000110_1=0;
q0000110_1=0;
m0000111_0=0;
q0000111_0=0;
m0000111_1=0;
q0000111_1=0;
m0001000_0=0;
q0001000_0=0;
m0001000_1=0;
q0001000_1=0;
m0001001_0=0;
q0001001_0=0;
m0001001_1=0;
q0001001_1=0;
m0001010_0=0;
q0001010_0=0;
m0001010_1=0;
q0001010_1=0;
m0001011_0=0;
q0001011_0=0;
m0001011_1=0;
q0001011_1=0;
m0001100_0=0;
q0001100_0=0;
m0001100_1=0;
q0001100_1=0;
m0001101_0=0;
q0001101_0=0;
m0001101_1=0;
q0001101_1=0;
m0001110_0=0;
q0001110_0=0;
m0001110_1=0;
q0001110_1=0;
m0001111_0=0;
q0001111_0=0;
m0001111_1=0;
q0001111_1=0;
m0010000_0=0;
q0010000_0=0;
m0010000_1=0;
q0010000_1=0;
m0010001_0=0;
q0010001_0=0;
m0010001_1=0;
q0010001_1=0;
m0010010_0=0;
q0010010_0=0;
m0010010_1=0;
q0010010_1=0;
m0010011_0=0;
q0010011_0=0;
m0010011_1=0;
q0010011_1=0;
m0010100_0=0;
q0010100_0=0;
m0010100_1=0;
q0010100_1=0;
m0010101_0=0;
q0010101_0=0;
m0010101_1=0;
q0010101_1=0;
m0010110_0=0;
q0010110_0=0;
m0010110_1=0;
q0010110_1=0;
m0010111_0=0;
q0010111_0=0;
m0010111_1=0;
q0010111_1=0;
m0011000_0=0;
q0011000_0=0;
m0011000_1=0;
q0011000_1=0;
m0011001_0=0;
q0011001_0=0;
m0011001_1=0;
q0011001_1=0;
m0011010_0=0;
q0011010_0=0;
m0011010_1=0;
q0011010_1=0;
m0011011_0=0;
q0011011_0=0;
m0011011_1=0;
q0011011_1=0;
m0011100_0=0;
q0011100_0=0;
m0011100_1=0;
q0011100_1=0;
m0011101_0=0;
q0011101_0=0;
m0011101_1=0;
q0011101_1=0;
m0011110_0=0;
q0011110_0=0;
m0011110_1=0;
q0011110_1=0;
m0011111_0=0;
q0011111_0=0;
m0011111_1=0;
q0011111_1=0;
m0100000_0=0;
q0100000_0=0;
m0100000_1=0;
q0100000_1=0;
m0100001_0=0;
q0100001_0=0;
m0100001_1=0;
q0100001_1=0;
m0100010_0=0;
q0100010_0=0;
m0100010_1=0;
q0100010_1=0;
m0100011_0=0;
q0100011_0=0;
m0100011_1=0;
q0100011_1=0;
m0100100_0=0;
q0100100_0=0;
m0100100_1=0;
q0100100_1=0;
m0100101_0=0;
q0100101_0=0;
m0100101_1=0;
q0100101_1=0;
m0100110_0=0;
q0100110_0=0;
m0100110_1=0;
q0100110_1=0;
m0100111_0=0;
q0100111_0=0;
m0100111_1=0;
q0100111_1=0;
m0101000_0=0;
q0101000_0=0;
m0101000_1=0;
q0101000_1=0;
m0101001_0=0;
q0101001_0=0;
m0101001_1=0;
q0101001_1=0;
m0101010_0=0;
q0101010_0=0;
m0101010_1=0;
q0101010_1=0;
m0101011_0=0;
q0101011_0=0;
m0101011_1=0;
q0101011_1=0;
m0101100_0=0;
q0101100_0=0;
m0101100_1=0;
q0101100_1=0;
m0101101_0=0;
q0101101_0=0;
m0101101_1=0;
q0101101_1=0;
m0101110_0=0;
q0101110_0=0;
m0101110_1=0;
q0101110_1=0;
m0101111_0=0;
q0101111_0=0;
m0101111_1=0;
q0101111_1=0;
m0110000_0=0;
q0110000_0=0;
m0110000_1=0;
q0110000_1=0;
m0110001_0=0;
q0110001_0=0;
m0110001_1=0;
q0110001_1=0;
m0110010_0=0;
q0110010_0=0;
m0110010_1=0;
q0110010_1=0;
m0110011_0=0;
q0110011_0=0;
m0110011_1=0;
q0110011_1=0;
m0110100_0=0;
q0110100_0=0;
m0110100_1=0;
q0110100_1=0;
m0110101_0=0;
q0110101_0=0;
m0110101_1=0;
q0110101_1=0;
m0110110_0=0;
q0110110_0=0;
m0110110_1=0;
q0110110_1=0;
m0110111_0=0;
q0110111_0=0;
m0110111_1=0;
q0110111_1=0;
m0111000_0=0;
q0111000_0=0;
m0111000_1=0;
q0111000_1=0;
m0111001_0=0;
q0111001_0=0;
m0111001_1=0;
q0111001_1=0;
m0111010_0=0;
q0111010_0=0;
m0111010_1=0;
q0111010_1=0;
m0111011_0=0;
q0111011_0=0;
m0111011_1=0;
q0111011_1=0;
m0111100_0=0;
q0111100_0=0;
m0111100_1=0;
q0111100_1=0;
m0111101_0=0;
q0111101_0=0;
m0111101_1=0;
q0111101_1=0;
m0111110_0=1;
q0111110_0=1;
m0111110_1=1;
q0111110_1=1;
m0111111_0=1;
q0111111_0=1;
m0111111_1=1;
q0111111_1=1;
m1000000_0=1;
q1000000_0=1;
m1000000_1=1;
q1000000_1=1;
m1000001_0=1;
q1000001_0=1;
m1000001_1=1;
q1000001_1=1;
m1000010_0=0;
q1000010_0=0;
m1000010_1=0;
q1000010_1=0;
m1000011_0=0;
q1000011_0=0;
m1000011_1=0;
q1000011_1=0;
m1000100_0=0;
q1000100_0=0;
m1000100_1=0;
q1000100_1=0;
m1000101_0=0;
q1000101_0=0;
m1000101_1=0;
q1000101_1=0;
m1000110_0=0;
q1000110_0=0;
m1000110_1=0;
q1000110_1=0;
m1000111_0=0;
q1000111_0=0;
m1000111_1=0;
q1000111_1=0;
m1001000_0=0;
q1001000_0=0;
m1001000_1=0;
q1001000_1=0;
m1001001_0=0;
q1001001_0=0;
m1001001_1=0;
q1001001_1=0;
m1001010_0=0;
q1001010_0=0;
m1001010_1=0;
q1001010_1=0;
m1001011_0=0;
q1001011_0=0;
m1001011_1=0;
q1001011_1=0;
m1001100_0=0;
q1001100_0=0;
m1001100_1=0;
q1001100_1=0;
m1001101_0=0;
q1001101_0=0;
m1001101_1=0;
q1001101_1=0;
m1001110_0=0;
q1001110_0=0;
m1001110_1=0;
q1001110_1=0;
m1001111_0=0;
q1001111_0=0;
m1001111_1=0;
q1001111_1=0;
m1010000_0=0;
q1010000_0=0;
m1010000_1=0;
q1010000_1=0;
m1010001_0=0;
q1010001_0=0;
m1010001_1=0;
q1010001_1=0;
m1010010_0=0;
q1010010_0=0;
m1010010_1=0;
q1010010_1=0;
m1010011_0=0;
q1010011_0=0;
m1010011_1=0;
q1010011_1=0;
m1010100_0=0;
q1010100_0=0;
m1010100_1=0;
q1010100_1=0;
m1010101_0=0;
q1010101_0=0;
m1010101_1=0;
q1010101_1=0;
m1010110_0=0;
q1010110_0=0;
m1010110_1=0;
q1010110_1=0;
m1010111_0=0;
q1010111_0=0;
m1010111_1=0;
q1010111_1=0;
m1011000_0=0;
q1011000_0=0;
m1011000_1=0;
q1011000_1=0;
m1011001_0=0;
q1011001_0=0;
m1011001_1=0;
q1011001_1=0;
m1011010_0=0;
q1011010_0=0;
m1011010_1=0;
q1011010_1=0;
m1011011_0=0;
q1011011_0=0;
m1011011_1=0;
q1011011_1=0;
m1011100_0=0;
q1011100_0=0;
m1011100_1=0;
q1011100_1=0;
m1011101_0=0;
q1011101_0=0;
m1011101_1=0;
q1011101_1=0;
m1011110_0=0;
q1011110_0=0;
m1011110_1=0;
q1011110_1=0;
m1011111_0=0;
q1011111_0=0;
m1011111_1=0;
q1011111_1=0;
m1100000_0=0;
q1100000_0=0;
m1100000_1=0;
q1100000_1=0;
m1100001_0=0;
q1100001_0=0;
m1100001_1=0;
q1100001_1=0;
m1100010_0=0;
q1100010_0=0;
m1100010_1=0;
q1100010_1=0;
m1100011_0=0;
q1100011_0=0;
m1100011_1=0;
q1100011_1=0;
m1100100_0=0;
q1100100_0=0;
m1100100_1=0;
q1100100_1=0;
m1100101_0=0;
q1100101_0=0;
m1100101_1=0;
q1100101_1=0;
m1100110_0=0;
q1100110_0=0;
m1100110_1=0;
q1100110_1=0;
m1100111_0=0;
q1100111_0=0;
m1100111_1=0;
q1100111_1=0;
m1101000_0=0;
q1101000_0=0;
m1101000_1=0;
q1101000_1=0;
m1101001_0=0;
q1101001_0=0;
m1101001_1=0;
q1101001_1=0;
m1101010_0=0;
q1101010_0=0;
m1101010_1=0;
q1101010_1=0;
m1101011_0=0;
q1101011_0=0;
m1101011_1=0;
q1101011_1=0;
m1101100_0=0;
q1101100_0=0;
m1101100_1=0;
q1101100_1=0;
m1101101_0=0;
q1101101_0=0;
m1101101_1=0;
q1101101_1=0;
m1101110_0=0;
q1101110_0=0;
m1101110_1=0;
q1101110_1=0;
m1101111_0=0;
q1101111_0=0;
m1101111_1=0;
q1101111_1=0;
m1110000_0=0;
q1110000_0=0;
m1110000_1=0;
q1110000_1=0;
m1110001_0=0;
q1110001_0=0;
m1110001_1=0;
q1110001_1=0;
m1110010_0=0;
q1110010_0=0;
m1110010_1=0;
q1110010_1=0;
m1110011_0=0;
q1110011_0=0;
m1110011_1=0;
q1110011_1=0;
m1110100_0=0;
q1110100_0=0;
m1110100_1=0;
q1110100_1=0;
m1110101_0=0;
q1110101_0=0;
m1110101_1=0;
q1110101_1=0;
m1110110_0=0;
q1110110_0=0;
m1110110_1=0;
q1110110_1=0;
m1110111_0=0;
q1110111_0=0;
m1110111_1=0;
q1110111_1=0;
m1111000_0=0;
q1111000_0=0;
m1111000_1=0;
q1111000_1=0;
m1111001_0=0;
q1111001_0=0;
m1111001_1=0;
q1111001_1=0;
m1111010_0=0;
q1111010_0=0;
m1111010_1=0;
q1111010_1=0;
m1111011_0=0;
q1111011_0=0;
m1111011_1=0;
q1111011_1=0;
m1111100_0=0;
q1111100_0=0;
m1111100_1=0;
q1111100_1=0;
m1111101_0=0;
q1111101_0=0;
m1111101_1=0;
q1111101_1=0;
m1111110_0=0;
q1111110_0=0;
m1111110_1=0;
q1111110_1=0;
m1111111_0=0;
q1111111_0=0;
m1111111_1=0;
q1111111_1=0;
m000000_0=1;
q000000_0=1;
m000000_1=1;
q000000_1=1;
m000001_0=1;
q000001_0=1;
m000001_1=1;
q000001_1=1;
m000010_0=0;
q000010_0=0;
m000010_1=0;
q000010_1=0;
m000011_0=0;
q000011_0=0;
m000011_1=0;
q000011_1=0;
m000100_0=0;
q000100_0=0;
m000100_1=0;
q000100_1=0;
m000101_0=0;
q000101_0=0;
m000101_1=0;
q000101_1=0;
m000110_0=0;
q000110_0=0;
m000110_1=0;
q000110_1=0;
m000111_0=0;
q000111_0=0;
m000111_1=0;
q000111_1=0;
m001000_0=0;
q001000_0=0;
m001000_1=0;
q001000_1=0;
m001001_0=0;
q001001_0=0;
m001001_1=0;
q001001_1=0;
m001010_0=0;
q001010_0=0;
m001010_1=0;
q001010_1=0;
m001011_0=0;
q001011_0=0;
m001011_1=0;
q001011_1=0;
m001100_0=0;
q001100_0=0;
m001100_1=0;
q001100_1=0;
m001101_0=0;
q001101_0=0;
m001101_1=0;
q001101_1=0;
m001110_0=0;
q001110_0=0;
m001110_1=0;
q001110_1=0;
m001111_0=0;
q001111_0=0;
m001111_1=0;
q001111_1=0;
m010000_0=0;
q010000_0=0;
m010000_1=0;
q010000_1=0;
m010001_0=0;
q010001_0=0;
m010001_1=0;
q010001_1=0;
m010010_0=0;
q010010_0=0;
m010010_1=0;
q010010_1=0;
m010011_0=0;
q010011_0=0;
m010011_1=0;
q010011_1=0;
m010100_0=0;
q010100_0=0;
m010100_1=0;
q010100_1=0;
m010101_0=0;
q010101_0=0;
m010101_1=0;
q010101_1=0;
m010110_0=0;
q010110_0=0;
m010110_1=0;
q010110_1=0;
m010111_0=0;
q010111_0=0;
m010111_1=0;
q010111_1=0;
m011000_0=0;
q011000_0=0;
m011000_1=0;
q011000_1=0;
m011001_0=0;
q011001_0=0;
m011001_1=0;
q011001_1=0;
m011010_0=0;
q011010_0=0;
m011010_1=0;
q011010_1=0;
m011011_0=0;
q011011_0=0;
m011011_1=0;
q011011_1=0;
m011100_0=0;
q011100_0=0;
m011100_1=0;
q011100_1=0;
m011101_0=0;
q011101_0=0;
m011101_1=0;
q011101_1=0;
m011110_0=1;
q011110_0=1;
m011110_1=1;
q011110_1=1;
m011111_0=1;
q011111_0=1;
m011111_1=1;
q011111_1=1;
m100000_0=1;
q100000_0=1;
m100000_1=1;
q100000_1=1;
m100001_0=1;
q100001_0=1;
m100001_1=1;
q100001_1=1;
m100010_0=0;
q100010_0=0;
m100010_1=0;
q100010_1=0;
m100011_0=0;
q100011_0=0;
m100011_1=0;
q100011_1=0;
m100100_0=0;
q100100_0=0;
m100100_1=0;
q100100_1=0;
m100101_0=0;
q100101_0=0;
m100101_1=0;
q100101_1=0;
m100110_0=0;
q100110_0=0;
m100110_1=0;
q100110_1=0;
m100111_0=0;
q100111_0=0;
m100111_1=0;
q100111_1=0;
m101000_0=0;
q101000_0=0;
m101000_1=0;
q101000_1=0;
m101001_0=0;
q101001_0=0;
m101001_1=0;
q101001_1=0;
m101010_0=0;
q101010_0=0;
m101010_1=0;
q101010_1=0;
m101011_0=0;
q101011_0=0;
m101011_1=0;
q101011_1=0;
m101100_0=0;
q101100_0=0;
m101100_1=0;
q101100_1=0;
m101101_0=0;
q101101_0=0;
m101101_1=0;
q101101_1=0;
m101110_0=0;
q101110_0=0;
m101110_1=0;
q101110_1=0;
m101111_0=0;
q101111_0=0;
m101111_1=0;
q101111_1=0;
m110000_0=0;
q110000_0=0;
m110000_1=0;
q110000_1=0;
m110001_0=0;
q110001_0=0;
m110001_1=0;
q110001_1=0;
m110010_0=0;
q110010_0=0;
m110010_1=0;
q110010_1=0;
m110011_0=0;
q110011_0=0;
m110011_1=0;
q110011_1=0;
m110100_0=0;
q110100_0=0;
m110100_1=0;
q110100_1=0;
m110101_0=0;
q110101_0=0;
m110101_1=0;
q110101_1=0;
m110110_0=0;
q110110_0=0;
m110110_1=0;
q110110_1=0;
m110111_0=0;
q110111_0=0;
m110111_1=0;
q110111_1=0;
m111000_0=0;
q111000_0=0;
m111000_1=0;
q111000_1=0;
m111001_0=0;
q111001_0=0;
m111001_1=0;
q111001_1=0;
m111010_0=0;
q111010_0=0;
m111010_1=0;
q111010_1=0;
m111011_0=0;
q111011_0=0;
m111011_1=0;
q111011_1=0;
m111100_0=0;
q111100_0=0;
m111100_1=0;
q111100_1=0;
m111101_0=0;
q111101_0=0;
m111101_1=0;
q111101_1=0;
m111110_0=1;
q111110_0=1;
m111110_1=1;
q111110_1=1;
m111111_0=1;
q111111_0=1;
m111111_1=1;
q111111_1=1;
m0061=1;
q0061=1;
m0062=1;
q0062=1;
m0063=1;
q0063=1;
m0064=1;
q0064=1;
m0065=1;
q0065=1;
m0066=1;
q0066=1;
m0067=1;
q0067=1;
m0068=1;
q0068=1;
m0069=1;
q0069=1;
m0070=1;
q0070=1;
m0071=1;
q0071=1;
m0072=1;
q0072=1;
m0073=1;
q0073=1;
m0074=1;
q0074=1;
m0075=1;
q0075=1;
m0076=1;
q0076=1;
m0077=1;
q0077=1;
m0078=1;
q0078=1;
m0079=1;
q0079=1;
m0080=1;
q0080=1;
m0081=0;
q0081=0;
m0082=0;
q0082=0;
m0083=0;
q0083=0;
m0084=0;
q0084=0;
m0085=0;
q0085=0;
m0086=0;
q0086=0;
m0087=0;
q0087=0;
m0088=0;
q0088=0;
m0089=0;
q0089=0;
m0090=0;
q0090=0;
m0121=1;
q0121=1;
m0122=1;
q0122=1;
m0123=1;
q0123=1;
m0124=1;
q0124=1;
m0125=1;
q0125=1;
m0126=1;
q0126=1;
m0127=1;
q0127=1;
m0128=1;
q0128=1;
m0129=1;
q0129=1;
m0130=1;
q0130=1;
m0131=1;
q0131=1;
m0132=1;
q0132=1;
m0133=1;
q0133=1;
m0134=1;
q0134=1;
m0135=1;
q0135=1;
m0136=1;
q0136=1;
m0137=1;
q0137=1;
m0138=1;
q0138=1;
m0139=1;
q0139=1;
m0140=1;
q0140=1;
m0141=1;
q0141=1;
m0142=1;
q0142=1;
m0143=1;
q0143=1;
m0144=0;
q0144=0;
m0145=0;
q0145=0;
m0146=0;
q0146=0;
m0147=0;
q0147=0;
m0148=0;
q0148=0;
m0149=0;
q0149=0;
m0150=0;
q0150=0;
m0181=1;
q0181=1;
m0182=1;
q0182=1;
m0183=1;
q0183=1;
m0184=1;
q0184=1;
m0185=1;
q0185=1;
m0186=1;
q0186=1;
m0187=1;
q0187=1;
m0188=1;
q0188=1;
m0189=1;
q0189=1;
m0190=1;
q0190=1;
m0191=1;
q0191=1;
m0192=1;
q0192=1;
m0193=1;
q0193=1;
m0194=1;
q0194=1;
m0195=1;
q0195=1;
m0196=1;
q0196=1;
m0197=1;
q0197=1;
m0198=1;
q0198=1;
m0199=1;
q0199=1;
m0200=1;
q0200=1;
m0201=0;
q0201=0;
m0202=0;
q0202=0;
m0203=0;
q0203=0;
m0204=0;
q0204=0;
m0205=0;
q0205=0;
m0206=0;
q0206=0;
m0207=0;
q0207=0;
m0208=0;
q0208=0;
m0209=0;
q0209=0;
m0210=0;
q0210=0;
m0241=1;
q0241=1;
m0242=1;
q0242=1;
m0243=1;
q0243=1;
m0244=1;
q0244=1;
m0245=1;
q0245=1;
m0246=1;
q0246=1;
m0247=1;
q0247=1;
m0248=1;
q0248=1;
m0249=1;
q0249=1;
m0250=1;
q0250=1;
m0251=1;
q0251=1;
m0252=1;
q0252=1;
m0253=1;
q0253=1;
m0254=1;
q0254=1;
m0255=1;
q0255=1;
m0256=1;
q0256=1;
m0257=1;
q0257=1;
m0258=1;
q0258=1;
m0259=1;
q0259=1;
m0260=1;
q0260=1;
m0261=0;
q0261=0;
m0262=0;
q0262=0;
m0263=0;
q0263=0;
m0264=0;
q0264=0;
m0265=0;
q0265=0;
m0266=0;
q0266=0;
m0267=0;
q0267=0;
m0268=0;
q0268=0;
m0269=0;
q0269=0;
m0270=0;
q0270=0;
m0301=1;
q0301=1;
m0302=1;
q0302=1;
m0303=1;
q0303=1;
m0304=1;
q0304=1;
m0305=1;
q0305=1;
m0306=1;
q0306=1;
m0307=1;
q0307=1;
m0308=1;
q0308=1;
m0309=0;
q0309=0;
m0310=0;
q0310=0;
m0311=1;
q0311=1;
m0312=1;
q0312=1;
m0313=0;
q0313=0;
m0314=1;
q0314=1;
m0315=0;
q0315=0;
m0316=0;
q0316=0;
m0317=1;
q0317=1;
m0318=0;
q0318=0;
m0319=0;
q0319=0;
m0320=0;
q0320=0;
m0321=1;
q0321=1;
m0322=1;
q0322=1;
m0323=0;
q0323=0;
m0324=0;
q0324=0;
m0325=1;
q0325=1;
m0326=0;
q0326=0;
m0327=0;
q0327=0;
m0328=0;
q0328=0;
m0329=0;
q0329=0;
m0330=0;
q0330=0;
m102_0=0;
q102_0=0;
m102_1=0;
q102_1=0;
m103_0=0;
q103_0=0;
m103_1=0;
q103_1=0;
m104_0=0;
q104_0=0;
m104_1=0;
q104_1=0;
m105_0=0;
q105_0=0;
m105_1=0;
q105_1=0;
m106_0=0;
q106_0=0;
m106_1=0;
q106_1=0;
m107_0=0;
q107_0=0;
m107_1=0;
q107_1=0;
m108_0=0;
q108_0=0;
m108_1=0;
q108_1=0;
m109_0=0;
q109_0=0;
m109_1=0;
q109_1=0;
m110_0=0;
q110_0=0;
m110_1=0;
q110_1=0;
m111_0=0;
q111_0=0;
m111_1=0;
q111_1=0;
m112_0=0;
q112_0=0;
m112_1=0;
q112_1=0;
m113_0=0;
q113_0=0;
m113_1=0;
q113_1=0;
m114_0=0;
q114_0=0;
m114_1=0;
q114_1=0;
m115_0=0;
q115_0=0;
m115_1=0;
q115_1=0;
m116_0=0;
q116_0=0;
m116_1=0;
q116_1=0;
m117_0=0;
q117_0=0;
m117_1=0;
q117_1=0;
m118_0=0;
q118_0=0;
m118_1=0;
q118_1=0;
m119_0=0;
q119_0=0;
m119_1=0;
q119_1=0;
m120_0=0;
q120_0=0;
m120_1=0;
q120_1=0;
m121_0=0;
q121_0=0;
m121_1=0;
q121_1=0;
m122_0=0;
q122_0=0;
m122_1=0;
q122_1=0;
m123_0=0;
q123_0=0;
m123_1=0;
q123_1=0;
m124_0=1;
q124_0=1;
m124_1=1;
q124_1=1;
m125_0=1;
q125_0=1;
m125_1=1;
q125_1=1;
m126_0=1;
q126_0=1;
m126_1=1;
q126_1=1;
m127_0=1;
q127_0=1;
m127_1=1;
q127_1=1;
m128_0=1;
q128_0=1;
m128_1=1;
q128_1=1;
m129_0=1;
q129_0=1;
m129_1=1;
q129_1=1;
m130_0=1;
q130_0=1;
m130_1=1;
q130_1=1;
m131_0=1;
q131_0=1;
m131_1=1;
q131_1=1;
m132_0=1;
q132_0=1;
m132_1=1;
q132_1=1;
m133_0=1;
q133_0=1;
m133_1=1;
q133_1=1;
m134_0=1;
q134_0=1;
m134_1=1;
q134_1=1;
m135_0=1;
q135_0=1;
m135_1=1;
q135_1=1;
m136_0=1;
q136_0=1;
m136_1=1;
q136_1=1;
m137_0=1;
q137_0=1;
m137_1=1;
q137_1=1;
m138_0=1;
q138_0=1;
m138_1=1;
q138_1=1;
m139_0=1;
q139_0=1;
m139_1=1;
q139_1=1;
m140_0=0;
q140_0=0;
m140_1=0;
q140_1=0;
m141_0=0;
q141_0=0;
m141_1=0;
q141_1=0;
m142_0=0;
q142_0=0;
m142_1=0;
q142_1=0;
m143_0=0;
q143_0=0;
m143_1=0;
q143_1=0;
m144_0=0;
q144_0=0;
m144_1=0;
q144_1=0;
m145_0=0;
q145_0=0;
m145_1=0;
q145_1=0;
m146_0=0;
q146_0=0;
m146_1=0;
q146_1=0;
m147_0=0;
q147_0=0;
m147_1=0;
q147_1=0;
m148_0=0;
q148_0=0;
m148_1=0;
q148_1=0;
m149_0=0;
q149_0=0;
m149_1=0;
q149_1=0;
m150_0=0;
q150_0=0;
m150_1=0;
q150_1=0;
m151_0=0;
q151_0=0;
m151_1=0;
q151_1=0;
m152_0=0;
q152_0=0;
m152_1=0;
q152_1=0;
m153_0=0;
q153_0=0;
m153_1=0;
q153_1=0;
m154_0=0;
q154_0=0;
m154_1=0;
q154_1=0;
m155_0=0;
q155_0=0;
m155_1=0;
q155_1=0;
m156_0=0;
q156_0=0;
m156_1=0;
q156_1=0;
m157_0=0;
q157_0=0;
m157_1=0;
q157_1=0;
m158_0=0;
q158_0=0;
m158_1=0;
q158_1=0;
m159_0=0;
q159_0=0;
m159_1=0;
q159_1=0;
m160_0=0;
q160_0=0;
m160_1=0;
q160_1=0;
m161_0=0;
q161_0=0;
m161_1=0;
q161_1=0;
m202_0=0;
q202_0=0;
m202_1=0;
q202_1=0;
m203_0=0;
q203_0=0;
m203_1=0;
q203_1=0;
m204_0=0;
q204_0=0;
m204_1=0;
q204_1=0;
m205_0=0;
q205_0=0;
m205_1=0;
q205_1=0;
m206_0=0;
q206_0=0;
m206_1=0;
q206_1=0;
m207_0=0;
q207_0=0;
m207_1=0;
q207_1=0;
m208_0=0;
q208_0=0;
m208_1=0;
q208_1=0;
m209_0=0;
q209_0=0;
m209_1=0;
q209_1=0;
m210_0=0;
q210_0=0;
m210_1=0;
q210_1=0;
m211_0=0;
q211_0=0;
m211_1=0;
q211_1=0;
m212_0=0;
q212_0=0;
m212_1=0;
q212_1=0;
m213_0=0;
q213_0=0;
m213_1=0;
q213_1=0;
m214_0=0;
q214_0=0;
m214_1=0;
q214_1=0;
m215_0=0;
q215_0=0;
m215_1=0;
q215_1=0;
m216_0=0;
q216_0=0;
m216_1=0;
q216_1=0;
m217_0=0;
q217_0=0;
m217_1=0;
q217_1=0;
m218_0=0;
q218_0=0;
m218_1=0;
q218_1=0;
m219_0=0;
q219_0=0;
m219_1=0;
q219_1=0;
m220_0=0;
q220_0=0;
m220_1=0;
q220_1=0;
m221_0=0;
q221_0=0;
m221_1=0;
q221_1=0;
m222_0=0;
q222_0=0;
m222_1=0;
q222_1=0;
m223_0=0;
q223_0=0;
m223_1=0;
q223_1=0;
m224_0=1;
q224_0=1;
m224_1=1;
q224_1=1;
m225_0=1;
q225_0=1;
m225_1=1;
q225_1=1;
m226_0=1;
q226_0=1;
m226_1=1;
q226_1=1;
m227_0=1;
q227_0=1;
m227_1=1;
q227_1=1;
m228_0=1;
q228_0=1;
m228_1=1;
q228_1=1;
m229_0=1;
q229_0=1;
m229_1=1;
q229_1=1;
m230_0=1;
q230_0=1;
m230_1=1;
q230_1=1;
m231_0=1;
q231_0=1;
m231_1=1;
q231_1=1;
m232_0=1;
q232_0=1;
m232_1=1;
q232_1=1;
m233_0=1;
q233_0=1;
m233_1=1;
q233_1=1;
m234_0=1;
q234_0=1;
m234_1=1;
q234_1=1;
m235_0=1;
q235_0=1;
m235_1=1;
q235_1=1;
m236_0=1;
q236_0=1;
m236_1=1;
q236_1=1;
m237_0=1;
q237_0=1;
m237_1=1;
q237_1=1;
m238_0=1;
q238_0=1;
m238_1=1;
q238_1=1;
m239_0=1;
q239_0=1;
m239_1=1;
q239_1=1;
m240_0=0;
q240_0=0;
m240_1=0;
q240_1=0;
m241_0=0;
q241_0=0;
m241_1=0;
q241_1=0;
m242_0=0;
q242_0=0;
m242_1=0;
q242_1=0;
m243_0=0;
q243_0=0;
m243_1=0;
q243_1=0;
m244_0=0;
q244_0=0;
m244_1=0;
q244_1=0;
m245_0=0;
q245_0=0;
m245_1=0;
q245_1=0;
m246_0=0;
q246_0=0;
m246_1=0;
q246_1=0;
m247_0=0;
q247_0=0;
m247_1=0;
q247_1=0;
m248_0=0;
q248_0=0;
m248_1=0;
q248_1=0;
m249_0=0;
q249_0=0;
m249_1=0;
q249_1=0;
m250_0=0;
q250_0=0;
m250_1=0;
q250_1=0;
m251_0=0;
q251_0=0;
m251_1=0;
q251_1=0;
m252_0=0;
q252_0=0;
m252_1=0;
q252_1=0;
m253_0=0;
q253_0=0;
m253_1=0;
q253_1=0;
m254_0=0;
q254_0=0;
m254_1=0;
q254_1=0;
m255_0=0;
q255_0=0;
m255_1=0;
q255_1=0;
m256_0=0;
q256_0=0;
m256_1=0;
q256_1=0;
m257_0=0;
q257_0=0;
m257_1=0;
q257_1=0;
m258_0=0;
q258_0=0;
m258_1=0;
q258_1=0;
m259_0=0;
q259_0=0;
m259_1=0;
q259_1=0;
m260_0=0;
q260_0=0;
m260_1=0;
q260_1=0;
m261_0=0;
q261_0=0;
m261_1=0;
q261_1=0;
m29_0=1;
q29_0=1;
m29_1=1;
q29_1=1;
m30_0=1;
q30_0=1;
m30_1=1;
q30_1=1;
m31_0=1;
q31_0=1;
m31_1=1;
q31_1=1;
m32_0=1;
q32_0=1;
m32_1=1;
q32_1=1;
m33_0=1;
q33_0=1;
m33_1=1;
q33_1=1;
m34_0=1;
q34_0=1;
m34_1=1;
q34_1=1;
m35_0=1;
q35_0=1;
m35_1=1;
q35_1=1;
m36_0=1;
q36_0=1;
m36_1=1;
q36_1=1;
m37_0=1;
q37_0=1;
m37_1=1;
q37_1=1;
m38_0=1;
q38_0=1;
m38_1=1;
q38_1=1;
m39_0=1;
q39_0=1;
m39_1=1;
q39_1=1;
m40_0=1;
q40_0=1;
m40_1=1;
q40_1=1;
m41_0=1;
q41_0=1;
m41_1=1;
q41_1=1;
m42_0=1;
q42_0=1;
m42_1=1;
q42_1=1;
m43_0=1;
q43_0=1;
m43_1=1;
q43_1=1;
m44_0=0;
q44_0=0;
m44_1=0;
q44_1=0;
m45_0=0;
q45_0=0;
m45_1=0;
q45_1=0;
m46_0=0;
q46_0=0;
m46_1=0;
q46_1=0;
m47_0=0;
q47_0=0;
m47_1=0;
q47_1=0;
m48_0=0;
q48_0=0;
m48_1=0;
q48_1=0;
m49_0=0;
q49_0=0;
m49_1=0;
q49_1=0;
m50_0=0;
q50_0=0;
m50_1=0;
q50_1=0;
end

endmodule
